module basic_PE(
  input         clock,
  input         reset,
  input  [7:0]  io_in_activate,
  input  [7:0]  io_in_weight,
  input  [15:0] io_in_psum,
  input         io_in_flow,
  input         io_in_shift,
  output [7:0]  io_out_activate,
  output [7:0]  io_out_weight,
  output [15:0] io_out_psum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] Activation_Reg; // @[basic_PE.scala 17:31]
  reg [7:0] Weight_Reg; // @[basic_PE.scala 18:27]
  reg [15:0] PSum_Reg; // @[basic_PE.scala 19:25]
  wire [15:0] _io_out_psum_T = Activation_Reg * Weight_Reg; // @[basic_PE.scala 47:33]
  assign io_out_activate = Activation_Reg; // @[basic_PE.scala 45:19]
  assign io_out_weight = Weight_Reg; // @[basic_PE.scala 46:17]
  assign io_out_psum = _io_out_psum_T + PSum_Reg; // @[basic_PE.scala 47:46]
  always @(posedge clock) begin
    if (reset) begin // @[basic_PE.scala 17:31]
      Activation_Reg <= 8'h0; // @[basic_PE.scala 17:31]
    end else if (io_in_flow) begin // @[basic_PE.scala 22:20]
      Activation_Reg <= io_in_activate; // @[basic_PE.scala 23:20]
    end
    if (reset) begin // @[basic_PE.scala 18:27]
      Weight_Reg <= 8'h0; // @[basic_PE.scala 18:27]
    end else if (io_in_shift) begin // @[basic_PE.scala 38:21]
      Weight_Reg <= io_in_weight; // @[basic_PE.scala 39:16]
    end
    if (reset) begin // @[basic_PE.scala 19:25]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 19:25]
    end else if (io_in_shift) begin // @[basic_PE.scala 29:21]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 30:14]
    end else if (io_in_flow) begin // @[basic_PE.scala 31:26]
      PSum_Reg <= io_in_psum; // @[basic_PE.scala 32:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Activation_Reg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  Weight_Reg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  PSum_Reg = _RAND_2[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Systolic_Array(
  input         clock,
  input         reset,
  input  [7:0]  io_activate_0,
  input  [7:0]  io_activate_1,
  input  [7:0]  io_activate_2,
  input  [7:0]  io_activate_3,
  input  [7:0]  io_activate_4,
  input  [7:0]  io_activate_5,
  input  [7:0]  io_activate_6,
  input  [7:0]  io_activate_7,
  input  [7:0]  io_activate_8,
  input  [7:0]  io_activate_9,
  input  [7:0]  io_activate_10,
  input  [7:0]  io_activate_11,
  input  [7:0]  io_activate_12,
  input  [7:0]  io_activate_13,
  input  [7:0]  io_activate_14,
  input  [7:0]  io_activate_15,
  input  [7:0]  io_weight_0,
  input  [7:0]  io_weight_1,
  input  [7:0]  io_weight_2,
  input  [7:0]  io_weight_3,
  input  [7:0]  io_weight_4,
  input  [7:0]  io_weight_5,
  input  [7:0]  io_weight_6,
  input  [7:0]  io_weight_7,
  input  [7:0]  io_weight_8,
  input  [7:0]  io_weight_9,
  input  [7:0]  io_weight_10,
  input  [7:0]  io_weight_11,
  input  [7:0]  io_weight_12,
  input  [7:0]  io_weight_13,
  input  [7:0]  io_weight_14,
  input  [7:0]  io_weight_15,
  input         io_flow,
  input         io_shift,
  output [15:0] io_psum_0,
  output [15:0] io_psum_1,
  output [15:0] io_psum_2,
  output [15:0] io_psum_3,
  output [15:0] io_psum_4,
  output [15:0] io_psum_5,
  output [15:0] io_psum_6,
  output [15:0] io_psum_7,
  output [15:0] io_psum_8,
  output [15:0] io_psum_9,
  output [15:0] io_psum_10,
  output [15:0] io_psum_11,
  output [15:0] io_psum_12,
  output [15:0] io_psum_13,
  output [15:0] io_psum_14,
  output [15:0] io_psum_15,
  output        io_valid_0,
  output        io_valid_1,
  output        io_valid_2,
  output        io_valid_3,
  output        io_valid_4,
  output        io_valid_5,
  output        io_valid_6,
  output        io_valid_7,
  output        io_valid_8,
  output        io_valid_9,
  output        io_valid_10,
  output        io_valid_11,
  output        io_valid_12,
  output        io_valid_13,
  output        io_valid_14,
  output        io_valid_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  PE_Array_0_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  reg [5:0] flow_counter; // @[Systolic_Array.scala 52:29]
  reg [15:0] valid_reg; // @[Systolic_Array.scala 53:26]
  wire [5:0] _flow_counter_T_1 = flow_counter + 6'h1; // @[Systolic_Array.scala 57:34]
  wire [15:0] _valid_reg_T_1 = {valid_reg[14:0],1'h1}; // @[Cat.scala 33:92]
  wire [15:0] _valid_reg_T_3 = {valid_reg[14:0],1'h0}; // @[Cat.scala 33:92]
  basic_PE PE_Array_0_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_0_clock),
    .reset(PE_Array_0_0_reset),
    .io_in_activate(PE_Array_0_0_io_in_activate),
    .io_in_weight(PE_Array_0_0_io_in_weight),
    .io_in_psum(PE_Array_0_0_io_in_psum),
    .io_in_flow(PE_Array_0_0_io_in_flow),
    .io_in_shift(PE_Array_0_0_io_in_shift),
    .io_out_activate(PE_Array_0_0_io_out_activate),
    .io_out_weight(PE_Array_0_0_io_out_weight),
    .io_out_psum(PE_Array_0_0_io_out_psum)
  );
  basic_PE PE_Array_0_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_1_clock),
    .reset(PE_Array_0_1_reset),
    .io_in_activate(PE_Array_0_1_io_in_activate),
    .io_in_weight(PE_Array_0_1_io_in_weight),
    .io_in_psum(PE_Array_0_1_io_in_psum),
    .io_in_flow(PE_Array_0_1_io_in_flow),
    .io_in_shift(PE_Array_0_1_io_in_shift),
    .io_out_activate(PE_Array_0_1_io_out_activate),
    .io_out_weight(PE_Array_0_1_io_out_weight),
    .io_out_psum(PE_Array_0_1_io_out_psum)
  );
  basic_PE PE_Array_0_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_2_clock),
    .reset(PE_Array_0_2_reset),
    .io_in_activate(PE_Array_0_2_io_in_activate),
    .io_in_weight(PE_Array_0_2_io_in_weight),
    .io_in_psum(PE_Array_0_2_io_in_psum),
    .io_in_flow(PE_Array_0_2_io_in_flow),
    .io_in_shift(PE_Array_0_2_io_in_shift),
    .io_out_activate(PE_Array_0_2_io_out_activate),
    .io_out_weight(PE_Array_0_2_io_out_weight),
    .io_out_psum(PE_Array_0_2_io_out_psum)
  );
  basic_PE PE_Array_0_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_3_clock),
    .reset(PE_Array_0_3_reset),
    .io_in_activate(PE_Array_0_3_io_in_activate),
    .io_in_weight(PE_Array_0_3_io_in_weight),
    .io_in_psum(PE_Array_0_3_io_in_psum),
    .io_in_flow(PE_Array_0_3_io_in_flow),
    .io_in_shift(PE_Array_0_3_io_in_shift),
    .io_out_activate(PE_Array_0_3_io_out_activate),
    .io_out_weight(PE_Array_0_3_io_out_weight),
    .io_out_psum(PE_Array_0_3_io_out_psum)
  );
  basic_PE PE_Array_0_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_4_clock),
    .reset(PE_Array_0_4_reset),
    .io_in_activate(PE_Array_0_4_io_in_activate),
    .io_in_weight(PE_Array_0_4_io_in_weight),
    .io_in_psum(PE_Array_0_4_io_in_psum),
    .io_in_flow(PE_Array_0_4_io_in_flow),
    .io_in_shift(PE_Array_0_4_io_in_shift),
    .io_out_activate(PE_Array_0_4_io_out_activate),
    .io_out_weight(PE_Array_0_4_io_out_weight),
    .io_out_psum(PE_Array_0_4_io_out_psum)
  );
  basic_PE PE_Array_0_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_5_clock),
    .reset(PE_Array_0_5_reset),
    .io_in_activate(PE_Array_0_5_io_in_activate),
    .io_in_weight(PE_Array_0_5_io_in_weight),
    .io_in_psum(PE_Array_0_5_io_in_psum),
    .io_in_flow(PE_Array_0_5_io_in_flow),
    .io_in_shift(PE_Array_0_5_io_in_shift),
    .io_out_activate(PE_Array_0_5_io_out_activate),
    .io_out_weight(PE_Array_0_5_io_out_weight),
    .io_out_psum(PE_Array_0_5_io_out_psum)
  );
  basic_PE PE_Array_0_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_6_clock),
    .reset(PE_Array_0_6_reset),
    .io_in_activate(PE_Array_0_6_io_in_activate),
    .io_in_weight(PE_Array_0_6_io_in_weight),
    .io_in_psum(PE_Array_0_6_io_in_psum),
    .io_in_flow(PE_Array_0_6_io_in_flow),
    .io_in_shift(PE_Array_0_6_io_in_shift),
    .io_out_activate(PE_Array_0_6_io_out_activate),
    .io_out_weight(PE_Array_0_6_io_out_weight),
    .io_out_psum(PE_Array_0_6_io_out_psum)
  );
  basic_PE PE_Array_0_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_7_clock),
    .reset(PE_Array_0_7_reset),
    .io_in_activate(PE_Array_0_7_io_in_activate),
    .io_in_weight(PE_Array_0_7_io_in_weight),
    .io_in_psum(PE_Array_0_7_io_in_psum),
    .io_in_flow(PE_Array_0_7_io_in_flow),
    .io_in_shift(PE_Array_0_7_io_in_shift),
    .io_out_activate(PE_Array_0_7_io_out_activate),
    .io_out_weight(PE_Array_0_7_io_out_weight),
    .io_out_psum(PE_Array_0_7_io_out_psum)
  );
  basic_PE PE_Array_0_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_8_clock),
    .reset(PE_Array_0_8_reset),
    .io_in_activate(PE_Array_0_8_io_in_activate),
    .io_in_weight(PE_Array_0_8_io_in_weight),
    .io_in_psum(PE_Array_0_8_io_in_psum),
    .io_in_flow(PE_Array_0_8_io_in_flow),
    .io_in_shift(PE_Array_0_8_io_in_shift),
    .io_out_activate(PE_Array_0_8_io_out_activate),
    .io_out_weight(PE_Array_0_8_io_out_weight),
    .io_out_psum(PE_Array_0_8_io_out_psum)
  );
  basic_PE PE_Array_0_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_9_clock),
    .reset(PE_Array_0_9_reset),
    .io_in_activate(PE_Array_0_9_io_in_activate),
    .io_in_weight(PE_Array_0_9_io_in_weight),
    .io_in_psum(PE_Array_0_9_io_in_psum),
    .io_in_flow(PE_Array_0_9_io_in_flow),
    .io_in_shift(PE_Array_0_9_io_in_shift),
    .io_out_activate(PE_Array_0_9_io_out_activate),
    .io_out_weight(PE_Array_0_9_io_out_weight),
    .io_out_psum(PE_Array_0_9_io_out_psum)
  );
  basic_PE PE_Array_0_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_10_clock),
    .reset(PE_Array_0_10_reset),
    .io_in_activate(PE_Array_0_10_io_in_activate),
    .io_in_weight(PE_Array_0_10_io_in_weight),
    .io_in_psum(PE_Array_0_10_io_in_psum),
    .io_in_flow(PE_Array_0_10_io_in_flow),
    .io_in_shift(PE_Array_0_10_io_in_shift),
    .io_out_activate(PE_Array_0_10_io_out_activate),
    .io_out_weight(PE_Array_0_10_io_out_weight),
    .io_out_psum(PE_Array_0_10_io_out_psum)
  );
  basic_PE PE_Array_0_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_11_clock),
    .reset(PE_Array_0_11_reset),
    .io_in_activate(PE_Array_0_11_io_in_activate),
    .io_in_weight(PE_Array_0_11_io_in_weight),
    .io_in_psum(PE_Array_0_11_io_in_psum),
    .io_in_flow(PE_Array_0_11_io_in_flow),
    .io_in_shift(PE_Array_0_11_io_in_shift),
    .io_out_activate(PE_Array_0_11_io_out_activate),
    .io_out_weight(PE_Array_0_11_io_out_weight),
    .io_out_psum(PE_Array_0_11_io_out_psum)
  );
  basic_PE PE_Array_0_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_12_clock),
    .reset(PE_Array_0_12_reset),
    .io_in_activate(PE_Array_0_12_io_in_activate),
    .io_in_weight(PE_Array_0_12_io_in_weight),
    .io_in_psum(PE_Array_0_12_io_in_psum),
    .io_in_flow(PE_Array_0_12_io_in_flow),
    .io_in_shift(PE_Array_0_12_io_in_shift),
    .io_out_activate(PE_Array_0_12_io_out_activate),
    .io_out_weight(PE_Array_0_12_io_out_weight),
    .io_out_psum(PE_Array_0_12_io_out_psum)
  );
  basic_PE PE_Array_0_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_13_clock),
    .reset(PE_Array_0_13_reset),
    .io_in_activate(PE_Array_0_13_io_in_activate),
    .io_in_weight(PE_Array_0_13_io_in_weight),
    .io_in_psum(PE_Array_0_13_io_in_psum),
    .io_in_flow(PE_Array_0_13_io_in_flow),
    .io_in_shift(PE_Array_0_13_io_in_shift),
    .io_out_activate(PE_Array_0_13_io_out_activate),
    .io_out_weight(PE_Array_0_13_io_out_weight),
    .io_out_psum(PE_Array_0_13_io_out_psum)
  );
  basic_PE PE_Array_0_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_14_clock),
    .reset(PE_Array_0_14_reset),
    .io_in_activate(PE_Array_0_14_io_in_activate),
    .io_in_weight(PE_Array_0_14_io_in_weight),
    .io_in_psum(PE_Array_0_14_io_in_psum),
    .io_in_flow(PE_Array_0_14_io_in_flow),
    .io_in_shift(PE_Array_0_14_io_in_shift),
    .io_out_activate(PE_Array_0_14_io_out_activate),
    .io_out_weight(PE_Array_0_14_io_out_weight),
    .io_out_psum(PE_Array_0_14_io_out_psum)
  );
  basic_PE PE_Array_0_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_15_clock),
    .reset(PE_Array_0_15_reset),
    .io_in_activate(PE_Array_0_15_io_in_activate),
    .io_in_weight(PE_Array_0_15_io_in_weight),
    .io_in_psum(PE_Array_0_15_io_in_psum),
    .io_in_flow(PE_Array_0_15_io_in_flow),
    .io_in_shift(PE_Array_0_15_io_in_shift),
    .io_out_activate(PE_Array_0_15_io_out_activate),
    .io_out_weight(PE_Array_0_15_io_out_weight),
    .io_out_psum(PE_Array_0_15_io_out_psum)
  );
  basic_PE PE_Array_1_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_0_clock),
    .reset(PE_Array_1_0_reset),
    .io_in_activate(PE_Array_1_0_io_in_activate),
    .io_in_weight(PE_Array_1_0_io_in_weight),
    .io_in_psum(PE_Array_1_0_io_in_psum),
    .io_in_flow(PE_Array_1_0_io_in_flow),
    .io_in_shift(PE_Array_1_0_io_in_shift),
    .io_out_activate(PE_Array_1_0_io_out_activate),
    .io_out_weight(PE_Array_1_0_io_out_weight),
    .io_out_psum(PE_Array_1_0_io_out_psum)
  );
  basic_PE PE_Array_1_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_1_clock),
    .reset(PE_Array_1_1_reset),
    .io_in_activate(PE_Array_1_1_io_in_activate),
    .io_in_weight(PE_Array_1_1_io_in_weight),
    .io_in_psum(PE_Array_1_1_io_in_psum),
    .io_in_flow(PE_Array_1_1_io_in_flow),
    .io_in_shift(PE_Array_1_1_io_in_shift),
    .io_out_activate(PE_Array_1_1_io_out_activate),
    .io_out_weight(PE_Array_1_1_io_out_weight),
    .io_out_psum(PE_Array_1_1_io_out_psum)
  );
  basic_PE PE_Array_1_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_2_clock),
    .reset(PE_Array_1_2_reset),
    .io_in_activate(PE_Array_1_2_io_in_activate),
    .io_in_weight(PE_Array_1_2_io_in_weight),
    .io_in_psum(PE_Array_1_2_io_in_psum),
    .io_in_flow(PE_Array_1_2_io_in_flow),
    .io_in_shift(PE_Array_1_2_io_in_shift),
    .io_out_activate(PE_Array_1_2_io_out_activate),
    .io_out_weight(PE_Array_1_2_io_out_weight),
    .io_out_psum(PE_Array_1_2_io_out_psum)
  );
  basic_PE PE_Array_1_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_3_clock),
    .reset(PE_Array_1_3_reset),
    .io_in_activate(PE_Array_1_3_io_in_activate),
    .io_in_weight(PE_Array_1_3_io_in_weight),
    .io_in_psum(PE_Array_1_3_io_in_psum),
    .io_in_flow(PE_Array_1_3_io_in_flow),
    .io_in_shift(PE_Array_1_3_io_in_shift),
    .io_out_activate(PE_Array_1_3_io_out_activate),
    .io_out_weight(PE_Array_1_3_io_out_weight),
    .io_out_psum(PE_Array_1_3_io_out_psum)
  );
  basic_PE PE_Array_1_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_4_clock),
    .reset(PE_Array_1_4_reset),
    .io_in_activate(PE_Array_1_4_io_in_activate),
    .io_in_weight(PE_Array_1_4_io_in_weight),
    .io_in_psum(PE_Array_1_4_io_in_psum),
    .io_in_flow(PE_Array_1_4_io_in_flow),
    .io_in_shift(PE_Array_1_4_io_in_shift),
    .io_out_activate(PE_Array_1_4_io_out_activate),
    .io_out_weight(PE_Array_1_4_io_out_weight),
    .io_out_psum(PE_Array_1_4_io_out_psum)
  );
  basic_PE PE_Array_1_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_5_clock),
    .reset(PE_Array_1_5_reset),
    .io_in_activate(PE_Array_1_5_io_in_activate),
    .io_in_weight(PE_Array_1_5_io_in_weight),
    .io_in_psum(PE_Array_1_5_io_in_psum),
    .io_in_flow(PE_Array_1_5_io_in_flow),
    .io_in_shift(PE_Array_1_5_io_in_shift),
    .io_out_activate(PE_Array_1_5_io_out_activate),
    .io_out_weight(PE_Array_1_5_io_out_weight),
    .io_out_psum(PE_Array_1_5_io_out_psum)
  );
  basic_PE PE_Array_1_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_6_clock),
    .reset(PE_Array_1_6_reset),
    .io_in_activate(PE_Array_1_6_io_in_activate),
    .io_in_weight(PE_Array_1_6_io_in_weight),
    .io_in_psum(PE_Array_1_6_io_in_psum),
    .io_in_flow(PE_Array_1_6_io_in_flow),
    .io_in_shift(PE_Array_1_6_io_in_shift),
    .io_out_activate(PE_Array_1_6_io_out_activate),
    .io_out_weight(PE_Array_1_6_io_out_weight),
    .io_out_psum(PE_Array_1_6_io_out_psum)
  );
  basic_PE PE_Array_1_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_7_clock),
    .reset(PE_Array_1_7_reset),
    .io_in_activate(PE_Array_1_7_io_in_activate),
    .io_in_weight(PE_Array_1_7_io_in_weight),
    .io_in_psum(PE_Array_1_7_io_in_psum),
    .io_in_flow(PE_Array_1_7_io_in_flow),
    .io_in_shift(PE_Array_1_7_io_in_shift),
    .io_out_activate(PE_Array_1_7_io_out_activate),
    .io_out_weight(PE_Array_1_7_io_out_weight),
    .io_out_psum(PE_Array_1_7_io_out_psum)
  );
  basic_PE PE_Array_1_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_8_clock),
    .reset(PE_Array_1_8_reset),
    .io_in_activate(PE_Array_1_8_io_in_activate),
    .io_in_weight(PE_Array_1_8_io_in_weight),
    .io_in_psum(PE_Array_1_8_io_in_psum),
    .io_in_flow(PE_Array_1_8_io_in_flow),
    .io_in_shift(PE_Array_1_8_io_in_shift),
    .io_out_activate(PE_Array_1_8_io_out_activate),
    .io_out_weight(PE_Array_1_8_io_out_weight),
    .io_out_psum(PE_Array_1_8_io_out_psum)
  );
  basic_PE PE_Array_1_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_9_clock),
    .reset(PE_Array_1_9_reset),
    .io_in_activate(PE_Array_1_9_io_in_activate),
    .io_in_weight(PE_Array_1_9_io_in_weight),
    .io_in_psum(PE_Array_1_9_io_in_psum),
    .io_in_flow(PE_Array_1_9_io_in_flow),
    .io_in_shift(PE_Array_1_9_io_in_shift),
    .io_out_activate(PE_Array_1_9_io_out_activate),
    .io_out_weight(PE_Array_1_9_io_out_weight),
    .io_out_psum(PE_Array_1_9_io_out_psum)
  );
  basic_PE PE_Array_1_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_10_clock),
    .reset(PE_Array_1_10_reset),
    .io_in_activate(PE_Array_1_10_io_in_activate),
    .io_in_weight(PE_Array_1_10_io_in_weight),
    .io_in_psum(PE_Array_1_10_io_in_psum),
    .io_in_flow(PE_Array_1_10_io_in_flow),
    .io_in_shift(PE_Array_1_10_io_in_shift),
    .io_out_activate(PE_Array_1_10_io_out_activate),
    .io_out_weight(PE_Array_1_10_io_out_weight),
    .io_out_psum(PE_Array_1_10_io_out_psum)
  );
  basic_PE PE_Array_1_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_11_clock),
    .reset(PE_Array_1_11_reset),
    .io_in_activate(PE_Array_1_11_io_in_activate),
    .io_in_weight(PE_Array_1_11_io_in_weight),
    .io_in_psum(PE_Array_1_11_io_in_psum),
    .io_in_flow(PE_Array_1_11_io_in_flow),
    .io_in_shift(PE_Array_1_11_io_in_shift),
    .io_out_activate(PE_Array_1_11_io_out_activate),
    .io_out_weight(PE_Array_1_11_io_out_weight),
    .io_out_psum(PE_Array_1_11_io_out_psum)
  );
  basic_PE PE_Array_1_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_12_clock),
    .reset(PE_Array_1_12_reset),
    .io_in_activate(PE_Array_1_12_io_in_activate),
    .io_in_weight(PE_Array_1_12_io_in_weight),
    .io_in_psum(PE_Array_1_12_io_in_psum),
    .io_in_flow(PE_Array_1_12_io_in_flow),
    .io_in_shift(PE_Array_1_12_io_in_shift),
    .io_out_activate(PE_Array_1_12_io_out_activate),
    .io_out_weight(PE_Array_1_12_io_out_weight),
    .io_out_psum(PE_Array_1_12_io_out_psum)
  );
  basic_PE PE_Array_1_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_13_clock),
    .reset(PE_Array_1_13_reset),
    .io_in_activate(PE_Array_1_13_io_in_activate),
    .io_in_weight(PE_Array_1_13_io_in_weight),
    .io_in_psum(PE_Array_1_13_io_in_psum),
    .io_in_flow(PE_Array_1_13_io_in_flow),
    .io_in_shift(PE_Array_1_13_io_in_shift),
    .io_out_activate(PE_Array_1_13_io_out_activate),
    .io_out_weight(PE_Array_1_13_io_out_weight),
    .io_out_psum(PE_Array_1_13_io_out_psum)
  );
  basic_PE PE_Array_1_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_14_clock),
    .reset(PE_Array_1_14_reset),
    .io_in_activate(PE_Array_1_14_io_in_activate),
    .io_in_weight(PE_Array_1_14_io_in_weight),
    .io_in_psum(PE_Array_1_14_io_in_psum),
    .io_in_flow(PE_Array_1_14_io_in_flow),
    .io_in_shift(PE_Array_1_14_io_in_shift),
    .io_out_activate(PE_Array_1_14_io_out_activate),
    .io_out_weight(PE_Array_1_14_io_out_weight),
    .io_out_psum(PE_Array_1_14_io_out_psum)
  );
  basic_PE PE_Array_1_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_15_clock),
    .reset(PE_Array_1_15_reset),
    .io_in_activate(PE_Array_1_15_io_in_activate),
    .io_in_weight(PE_Array_1_15_io_in_weight),
    .io_in_psum(PE_Array_1_15_io_in_psum),
    .io_in_flow(PE_Array_1_15_io_in_flow),
    .io_in_shift(PE_Array_1_15_io_in_shift),
    .io_out_activate(PE_Array_1_15_io_out_activate),
    .io_out_weight(PE_Array_1_15_io_out_weight),
    .io_out_psum(PE_Array_1_15_io_out_psum)
  );
  basic_PE PE_Array_2_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_0_clock),
    .reset(PE_Array_2_0_reset),
    .io_in_activate(PE_Array_2_0_io_in_activate),
    .io_in_weight(PE_Array_2_0_io_in_weight),
    .io_in_psum(PE_Array_2_0_io_in_psum),
    .io_in_flow(PE_Array_2_0_io_in_flow),
    .io_in_shift(PE_Array_2_0_io_in_shift),
    .io_out_activate(PE_Array_2_0_io_out_activate),
    .io_out_weight(PE_Array_2_0_io_out_weight),
    .io_out_psum(PE_Array_2_0_io_out_psum)
  );
  basic_PE PE_Array_2_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_1_clock),
    .reset(PE_Array_2_1_reset),
    .io_in_activate(PE_Array_2_1_io_in_activate),
    .io_in_weight(PE_Array_2_1_io_in_weight),
    .io_in_psum(PE_Array_2_1_io_in_psum),
    .io_in_flow(PE_Array_2_1_io_in_flow),
    .io_in_shift(PE_Array_2_1_io_in_shift),
    .io_out_activate(PE_Array_2_1_io_out_activate),
    .io_out_weight(PE_Array_2_1_io_out_weight),
    .io_out_psum(PE_Array_2_1_io_out_psum)
  );
  basic_PE PE_Array_2_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_2_clock),
    .reset(PE_Array_2_2_reset),
    .io_in_activate(PE_Array_2_2_io_in_activate),
    .io_in_weight(PE_Array_2_2_io_in_weight),
    .io_in_psum(PE_Array_2_2_io_in_psum),
    .io_in_flow(PE_Array_2_2_io_in_flow),
    .io_in_shift(PE_Array_2_2_io_in_shift),
    .io_out_activate(PE_Array_2_2_io_out_activate),
    .io_out_weight(PE_Array_2_2_io_out_weight),
    .io_out_psum(PE_Array_2_2_io_out_psum)
  );
  basic_PE PE_Array_2_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_3_clock),
    .reset(PE_Array_2_3_reset),
    .io_in_activate(PE_Array_2_3_io_in_activate),
    .io_in_weight(PE_Array_2_3_io_in_weight),
    .io_in_psum(PE_Array_2_3_io_in_psum),
    .io_in_flow(PE_Array_2_3_io_in_flow),
    .io_in_shift(PE_Array_2_3_io_in_shift),
    .io_out_activate(PE_Array_2_3_io_out_activate),
    .io_out_weight(PE_Array_2_3_io_out_weight),
    .io_out_psum(PE_Array_2_3_io_out_psum)
  );
  basic_PE PE_Array_2_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_4_clock),
    .reset(PE_Array_2_4_reset),
    .io_in_activate(PE_Array_2_4_io_in_activate),
    .io_in_weight(PE_Array_2_4_io_in_weight),
    .io_in_psum(PE_Array_2_4_io_in_psum),
    .io_in_flow(PE_Array_2_4_io_in_flow),
    .io_in_shift(PE_Array_2_4_io_in_shift),
    .io_out_activate(PE_Array_2_4_io_out_activate),
    .io_out_weight(PE_Array_2_4_io_out_weight),
    .io_out_psum(PE_Array_2_4_io_out_psum)
  );
  basic_PE PE_Array_2_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_5_clock),
    .reset(PE_Array_2_5_reset),
    .io_in_activate(PE_Array_2_5_io_in_activate),
    .io_in_weight(PE_Array_2_5_io_in_weight),
    .io_in_psum(PE_Array_2_5_io_in_psum),
    .io_in_flow(PE_Array_2_5_io_in_flow),
    .io_in_shift(PE_Array_2_5_io_in_shift),
    .io_out_activate(PE_Array_2_5_io_out_activate),
    .io_out_weight(PE_Array_2_5_io_out_weight),
    .io_out_psum(PE_Array_2_5_io_out_psum)
  );
  basic_PE PE_Array_2_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_6_clock),
    .reset(PE_Array_2_6_reset),
    .io_in_activate(PE_Array_2_6_io_in_activate),
    .io_in_weight(PE_Array_2_6_io_in_weight),
    .io_in_psum(PE_Array_2_6_io_in_psum),
    .io_in_flow(PE_Array_2_6_io_in_flow),
    .io_in_shift(PE_Array_2_6_io_in_shift),
    .io_out_activate(PE_Array_2_6_io_out_activate),
    .io_out_weight(PE_Array_2_6_io_out_weight),
    .io_out_psum(PE_Array_2_6_io_out_psum)
  );
  basic_PE PE_Array_2_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_7_clock),
    .reset(PE_Array_2_7_reset),
    .io_in_activate(PE_Array_2_7_io_in_activate),
    .io_in_weight(PE_Array_2_7_io_in_weight),
    .io_in_psum(PE_Array_2_7_io_in_psum),
    .io_in_flow(PE_Array_2_7_io_in_flow),
    .io_in_shift(PE_Array_2_7_io_in_shift),
    .io_out_activate(PE_Array_2_7_io_out_activate),
    .io_out_weight(PE_Array_2_7_io_out_weight),
    .io_out_psum(PE_Array_2_7_io_out_psum)
  );
  basic_PE PE_Array_2_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_8_clock),
    .reset(PE_Array_2_8_reset),
    .io_in_activate(PE_Array_2_8_io_in_activate),
    .io_in_weight(PE_Array_2_8_io_in_weight),
    .io_in_psum(PE_Array_2_8_io_in_psum),
    .io_in_flow(PE_Array_2_8_io_in_flow),
    .io_in_shift(PE_Array_2_8_io_in_shift),
    .io_out_activate(PE_Array_2_8_io_out_activate),
    .io_out_weight(PE_Array_2_8_io_out_weight),
    .io_out_psum(PE_Array_2_8_io_out_psum)
  );
  basic_PE PE_Array_2_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_9_clock),
    .reset(PE_Array_2_9_reset),
    .io_in_activate(PE_Array_2_9_io_in_activate),
    .io_in_weight(PE_Array_2_9_io_in_weight),
    .io_in_psum(PE_Array_2_9_io_in_psum),
    .io_in_flow(PE_Array_2_9_io_in_flow),
    .io_in_shift(PE_Array_2_9_io_in_shift),
    .io_out_activate(PE_Array_2_9_io_out_activate),
    .io_out_weight(PE_Array_2_9_io_out_weight),
    .io_out_psum(PE_Array_2_9_io_out_psum)
  );
  basic_PE PE_Array_2_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_10_clock),
    .reset(PE_Array_2_10_reset),
    .io_in_activate(PE_Array_2_10_io_in_activate),
    .io_in_weight(PE_Array_2_10_io_in_weight),
    .io_in_psum(PE_Array_2_10_io_in_psum),
    .io_in_flow(PE_Array_2_10_io_in_flow),
    .io_in_shift(PE_Array_2_10_io_in_shift),
    .io_out_activate(PE_Array_2_10_io_out_activate),
    .io_out_weight(PE_Array_2_10_io_out_weight),
    .io_out_psum(PE_Array_2_10_io_out_psum)
  );
  basic_PE PE_Array_2_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_11_clock),
    .reset(PE_Array_2_11_reset),
    .io_in_activate(PE_Array_2_11_io_in_activate),
    .io_in_weight(PE_Array_2_11_io_in_weight),
    .io_in_psum(PE_Array_2_11_io_in_psum),
    .io_in_flow(PE_Array_2_11_io_in_flow),
    .io_in_shift(PE_Array_2_11_io_in_shift),
    .io_out_activate(PE_Array_2_11_io_out_activate),
    .io_out_weight(PE_Array_2_11_io_out_weight),
    .io_out_psum(PE_Array_2_11_io_out_psum)
  );
  basic_PE PE_Array_2_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_12_clock),
    .reset(PE_Array_2_12_reset),
    .io_in_activate(PE_Array_2_12_io_in_activate),
    .io_in_weight(PE_Array_2_12_io_in_weight),
    .io_in_psum(PE_Array_2_12_io_in_psum),
    .io_in_flow(PE_Array_2_12_io_in_flow),
    .io_in_shift(PE_Array_2_12_io_in_shift),
    .io_out_activate(PE_Array_2_12_io_out_activate),
    .io_out_weight(PE_Array_2_12_io_out_weight),
    .io_out_psum(PE_Array_2_12_io_out_psum)
  );
  basic_PE PE_Array_2_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_13_clock),
    .reset(PE_Array_2_13_reset),
    .io_in_activate(PE_Array_2_13_io_in_activate),
    .io_in_weight(PE_Array_2_13_io_in_weight),
    .io_in_psum(PE_Array_2_13_io_in_psum),
    .io_in_flow(PE_Array_2_13_io_in_flow),
    .io_in_shift(PE_Array_2_13_io_in_shift),
    .io_out_activate(PE_Array_2_13_io_out_activate),
    .io_out_weight(PE_Array_2_13_io_out_weight),
    .io_out_psum(PE_Array_2_13_io_out_psum)
  );
  basic_PE PE_Array_2_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_14_clock),
    .reset(PE_Array_2_14_reset),
    .io_in_activate(PE_Array_2_14_io_in_activate),
    .io_in_weight(PE_Array_2_14_io_in_weight),
    .io_in_psum(PE_Array_2_14_io_in_psum),
    .io_in_flow(PE_Array_2_14_io_in_flow),
    .io_in_shift(PE_Array_2_14_io_in_shift),
    .io_out_activate(PE_Array_2_14_io_out_activate),
    .io_out_weight(PE_Array_2_14_io_out_weight),
    .io_out_psum(PE_Array_2_14_io_out_psum)
  );
  basic_PE PE_Array_2_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_15_clock),
    .reset(PE_Array_2_15_reset),
    .io_in_activate(PE_Array_2_15_io_in_activate),
    .io_in_weight(PE_Array_2_15_io_in_weight),
    .io_in_psum(PE_Array_2_15_io_in_psum),
    .io_in_flow(PE_Array_2_15_io_in_flow),
    .io_in_shift(PE_Array_2_15_io_in_shift),
    .io_out_activate(PE_Array_2_15_io_out_activate),
    .io_out_weight(PE_Array_2_15_io_out_weight),
    .io_out_psum(PE_Array_2_15_io_out_psum)
  );
  basic_PE PE_Array_3_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_0_clock),
    .reset(PE_Array_3_0_reset),
    .io_in_activate(PE_Array_3_0_io_in_activate),
    .io_in_weight(PE_Array_3_0_io_in_weight),
    .io_in_psum(PE_Array_3_0_io_in_psum),
    .io_in_flow(PE_Array_3_0_io_in_flow),
    .io_in_shift(PE_Array_3_0_io_in_shift),
    .io_out_activate(PE_Array_3_0_io_out_activate),
    .io_out_weight(PE_Array_3_0_io_out_weight),
    .io_out_psum(PE_Array_3_0_io_out_psum)
  );
  basic_PE PE_Array_3_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_1_clock),
    .reset(PE_Array_3_1_reset),
    .io_in_activate(PE_Array_3_1_io_in_activate),
    .io_in_weight(PE_Array_3_1_io_in_weight),
    .io_in_psum(PE_Array_3_1_io_in_psum),
    .io_in_flow(PE_Array_3_1_io_in_flow),
    .io_in_shift(PE_Array_3_1_io_in_shift),
    .io_out_activate(PE_Array_3_1_io_out_activate),
    .io_out_weight(PE_Array_3_1_io_out_weight),
    .io_out_psum(PE_Array_3_1_io_out_psum)
  );
  basic_PE PE_Array_3_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_2_clock),
    .reset(PE_Array_3_2_reset),
    .io_in_activate(PE_Array_3_2_io_in_activate),
    .io_in_weight(PE_Array_3_2_io_in_weight),
    .io_in_psum(PE_Array_3_2_io_in_psum),
    .io_in_flow(PE_Array_3_2_io_in_flow),
    .io_in_shift(PE_Array_3_2_io_in_shift),
    .io_out_activate(PE_Array_3_2_io_out_activate),
    .io_out_weight(PE_Array_3_2_io_out_weight),
    .io_out_psum(PE_Array_3_2_io_out_psum)
  );
  basic_PE PE_Array_3_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_3_clock),
    .reset(PE_Array_3_3_reset),
    .io_in_activate(PE_Array_3_3_io_in_activate),
    .io_in_weight(PE_Array_3_3_io_in_weight),
    .io_in_psum(PE_Array_3_3_io_in_psum),
    .io_in_flow(PE_Array_3_3_io_in_flow),
    .io_in_shift(PE_Array_3_3_io_in_shift),
    .io_out_activate(PE_Array_3_3_io_out_activate),
    .io_out_weight(PE_Array_3_3_io_out_weight),
    .io_out_psum(PE_Array_3_3_io_out_psum)
  );
  basic_PE PE_Array_3_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_4_clock),
    .reset(PE_Array_3_4_reset),
    .io_in_activate(PE_Array_3_4_io_in_activate),
    .io_in_weight(PE_Array_3_4_io_in_weight),
    .io_in_psum(PE_Array_3_4_io_in_psum),
    .io_in_flow(PE_Array_3_4_io_in_flow),
    .io_in_shift(PE_Array_3_4_io_in_shift),
    .io_out_activate(PE_Array_3_4_io_out_activate),
    .io_out_weight(PE_Array_3_4_io_out_weight),
    .io_out_psum(PE_Array_3_4_io_out_psum)
  );
  basic_PE PE_Array_3_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_5_clock),
    .reset(PE_Array_3_5_reset),
    .io_in_activate(PE_Array_3_5_io_in_activate),
    .io_in_weight(PE_Array_3_5_io_in_weight),
    .io_in_psum(PE_Array_3_5_io_in_psum),
    .io_in_flow(PE_Array_3_5_io_in_flow),
    .io_in_shift(PE_Array_3_5_io_in_shift),
    .io_out_activate(PE_Array_3_5_io_out_activate),
    .io_out_weight(PE_Array_3_5_io_out_weight),
    .io_out_psum(PE_Array_3_5_io_out_psum)
  );
  basic_PE PE_Array_3_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_6_clock),
    .reset(PE_Array_3_6_reset),
    .io_in_activate(PE_Array_3_6_io_in_activate),
    .io_in_weight(PE_Array_3_6_io_in_weight),
    .io_in_psum(PE_Array_3_6_io_in_psum),
    .io_in_flow(PE_Array_3_6_io_in_flow),
    .io_in_shift(PE_Array_3_6_io_in_shift),
    .io_out_activate(PE_Array_3_6_io_out_activate),
    .io_out_weight(PE_Array_3_6_io_out_weight),
    .io_out_psum(PE_Array_3_6_io_out_psum)
  );
  basic_PE PE_Array_3_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_7_clock),
    .reset(PE_Array_3_7_reset),
    .io_in_activate(PE_Array_3_7_io_in_activate),
    .io_in_weight(PE_Array_3_7_io_in_weight),
    .io_in_psum(PE_Array_3_7_io_in_psum),
    .io_in_flow(PE_Array_3_7_io_in_flow),
    .io_in_shift(PE_Array_3_7_io_in_shift),
    .io_out_activate(PE_Array_3_7_io_out_activate),
    .io_out_weight(PE_Array_3_7_io_out_weight),
    .io_out_psum(PE_Array_3_7_io_out_psum)
  );
  basic_PE PE_Array_3_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_8_clock),
    .reset(PE_Array_3_8_reset),
    .io_in_activate(PE_Array_3_8_io_in_activate),
    .io_in_weight(PE_Array_3_8_io_in_weight),
    .io_in_psum(PE_Array_3_8_io_in_psum),
    .io_in_flow(PE_Array_3_8_io_in_flow),
    .io_in_shift(PE_Array_3_8_io_in_shift),
    .io_out_activate(PE_Array_3_8_io_out_activate),
    .io_out_weight(PE_Array_3_8_io_out_weight),
    .io_out_psum(PE_Array_3_8_io_out_psum)
  );
  basic_PE PE_Array_3_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_9_clock),
    .reset(PE_Array_3_9_reset),
    .io_in_activate(PE_Array_3_9_io_in_activate),
    .io_in_weight(PE_Array_3_9_io_in_weight),
    .io_in_psum(PE_Array_3_9_io_in_psum),
    .io_in_flow(PE_Array_3_9_io_in_flow),
    .io_in_shift(PE_Array_3_9_io_in_shift),
    .io_out_activate(PE_Array_3_9_io_out_activate),
    .io_out_weight(PE_Array_3_9_io_out_weight),
    .io_out_psum(PE_Array_3_9_io_out_psum)
  );
  basic_PE PE_Array_3_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_10_clock),
    .reset(PE_Array_3_10_reset),
    .io_in_activate(PE_Array_3_10_io_in_activate),
    .io_in_weight(PE_Array_3_10_io_in_weight),
    .io_in_psum(PE_Array_3_10_io_in_psum),
    .io_in_flow(PE_Array_3_10_io_in_flow),
    .io_in_shift(PE_Array_3_10_io_in_shift),
    .io_out_activate(PE_Array_3_10_io_out_activate),
    .io_out_weight(PE_Array_3_10_io_out_weight),
    .io_out_psum(PE_Array_3_10_io_out_psum)
  );
  basic_PE PE_Array_3_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_11_clock),
    .reset(PE_Array_3_11_reset),
    .io_in_activate(PE_Array_3_11_io_in_activate),
    .io_in_weight(PE_Array_3_11_io_in_weight),
    .io_in_psum(PE_Array_3_11_io_in_psum),
    .io_in_flow(PE_Array_3_11_io_in_flow),
    .io_in_shift(PE_Array_3_11_io_in_shift),
    .io_out_activate(PE_Array_3_11_io_out_activate),
    .io_out_weight(PE_Array_3_11_io_out_weight),
    .io_out_psum(PE_Array_3_11_io_out_psum)
  );
  basic_PE PE_Array_3_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_12_clock),
    .reset(PE_Array_3_12_reset),
    .io_in_activate(PE_Array_3_12_io_in_activate),
    .io_in_weight(PE_Array_3_12_io_in_weight),
    .io_in_psum(PE_Array_3_12_io_in_psum),
    .io_in_flow(PE_Array_3_12_io_in_flow),
    .io_in_shift(PE_Array_3_12_io_in_shift),
    .io_out_activate(PE_Array_3_12_io_out_activate),
    .io_out_weight(PE_Array_3_12_io_out_weight),
    .io_out_psum(PE_Array_3_12_io_out_psum)
  );
  basic_PE PE_Array_3_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_13_clock),
    .reset(PE_Array_3_13_reset),
    .io_in_activate(PE_Array_3_13_io_in_activate),
    .io_in_weight(PE_Array_3_13_io_in_weight),
    .io_in_psum(PE_Array_3_13_io_in_psum),
    .io_in_flow(PE_Array_3_13_io_in_flow),
    .io_in_shift(PE_Array_3_13_io_in_shift),
    .io_out_activate(PE_Array_3_13_io_out_activate),
    .io_out_weight(PE_Array_3_13_io_out_weight),
    .io_out_psum(PE_Array_3_13_io_out_psum)
  );
  basic_PE PE_Array_3_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_14_clock),
    .reset(PE_Array_3_14_reset),
    .io_in_activate(PE_Array_3_14_io_in_activate),
    .io_in_weight(PE_Array_3_14_io_in_weight),
    .io_in_psum(PE_Array_3_14_io_in_psum),
    .io_in_flow(PE_Array_3_14_io_in_flow),
    .io_in_shift(PE_Array_3_14_io_in_shift),
    .io_out_activate(PE_Array_3_14_io_out_activate),
    .io_out_weight(PE_Array_3_14_io_out_weight),
    .io_out_psum(PE_Array_3_14_io_out_psum)
  );
  basic_PE PE_Array_3_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_15_clock),
    .reset(PE_Array_3_15_reset),
    .io_in_activate(PE_Array_3_15_io_in_activate),
    .io_in_weight(PE_Array_3_15_io_in_weight),
    .io_in_psum(PE_Array_3_15_io_in_psum),
    .io_in_flow(PE_Array_3_15_io_in_flow),
    .io_in_shift(PE_Array_3_15_io_in_shift),
    .io_out_activate(PE_Array_3_15_io_out_activate),
    .io_out_weight(PE_Array_3_15_io_out_weight),
    .io_out_psum(PE_Array_3_15_io_out_psum)
  );
  basic_PE PE_Array_4_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_0_clock),
    .reset(PE_Array_4_0_reset),
    .io_in_activate(PE_Array_4_0_io_in_activate),
    .io_in_weight(PE_Array_4_0_io_in_weight),
    .io_in_psum(PE_Array_4_0_io_in_psum),
    .io_in_flow(PE_Array_4_0_io_in_flow),
    .io_in_shift(PE_Array_4_0_io_in_shift),
    .io_out_activate(PE_Array_4_0_io_out_activate),
    .io_out_weight(PE_Array_4_0_io_out_weight),
    .io_out_psum(PE_Array_4_0_io_out_psum)
  );
  basic_PE PE_Array_4_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_1_clock),
    .reset(PE_Array_4_1_reset),
    .io_in_activate(PE_Array_4_1_io_in_activate),
    .io_in_weight(PE_Array_4_1_io_in_weight),
    .io_in_psum(PE_Array_4_1_io_in_psum),
    .io_in_flow(PE_Array_4_1_io_in_flow),
    .io_in_shift(PE_Array_4_1_io_in_shift),
    .io_out_activate(PE_Array_4_1_io_out_activate),
    .io_out_weight(PE_Array_4_1_io_out_weight),
    .io_out_psum(PE_Array_4_1_io_out_psum)
  );
  basic_PE PE_Array_4_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_2_clock),
    .reset(PE_Array_4_2_reset),
    .io_in_activate(PE_Array_4_2_io_in_activate),
    .io_in_weight(PE_Array_4_2_io_in_weight),
    .io_in_psum(PE_Array_4_2_io_in_psum),
    .io_in_flow(PE_Array_4_2_io_in_flow),
    .io_in_shift(PE_Array_4_2_io_in_shift),
    .io_out_activate(PE_Array_4_2_io_out_activate),
    .io_out_weight(PE_Array_4_2_io_out_weight),
    .io_out_psum(PE_Array_4_2_io_out_psum)
  );
  basic_PE PE_Array_4_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_3_clock),
    .reset(PE_Array_4_3_reset),
    .io_in_activate(PE_Array_4_3_io_in_activate),
    .io_in_weight(PE_Array_4_3_io_in_weight),
    .io_in_psum(PE_Array_4_3_io_in_psum),
    .io_in_flow(PE_Array_4_3_io_in_flow),
    .io_in_shift(PE_Array_4_3_io_in_shift),
    .io_out_activate(PE_Array_4_3_io_out_activate),
    .io_out_weight(PE_Array_4_3_io_out_weight),
    .io_out_psum(PE_Array_4_3_io_out_psum)
  );
  basic_PE PE_Array_4_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_4_clock),
    .reset(PE_Array_4_4_reset),
    .io_in_activate(PE_Array_4_4_io_in_activate),
    .io_in_weight(PE_Array_4_4_io_in_weight),
    .io_in_psum(PE_Array_4_4_io_in_psum),
    .io_in_flow(PE_Array_4_4_io_in_flow),
    .io_in_shift(PE_Array_4_4_io_in_shift),
    .io_out_activate(PE_Array_4_4_io_out_activate),
    .io_out_weight(PE_Array_4_4_io_out_weight),
    .io_out_psum(PE_Array_4_4_io_out_psum)
  );
  basic_PE PE_Array_4_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_5_clock),
    .reset(PE_Array_4_5_reset),
    .io_in_activate(PE_Array_4_5_io_in_activate),
    .io_in_weight(PE_Array_4_5_io_in_weight),
    .io_in_psum(PE_Array_4_5_io_in_psum),
    .io_in_flow(PE_Array_4_5_io_in_flow),
    .io_in_shift(PE_Array_4_5_io_in_shift),
    .io_out_activate(PE_Array_4_5_io_out_activate),
    .io_out_weight(PE_Array_4_5_io_out_weight),
    .io_out_psum(PE_Array_4_5_io_out_psum)
  );
  basic_PE PE_Array_4_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_6_clock),
    .reset(PE_Array_4_6_reset),
    .io_in_activate(PE_Array_4_6_io_in_activate),
    .io_in_weight(PE_Array_4_6_io_in_weight),
    .io_in_psum(PE_Array_4_6_io_in_psum),
    .io_in_flow(PE_Array_4_6_io_in_flow),
    .io_in_shift(PE_Array_4_6_io_in_shift),
    .io_out_activate(PE_Array_4_6_io_out_activate),
    .io_out_weight(PE_Array_4_6_io_out_weight),
    .io_out_psum(PE_Array_4_6_io_out_psum)
  );
  basic_PE PE_Array_4_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_7_clock),
    .reset(PE_Array_4_7_reset),
    .io_in_activate(PE_Array_4_7_io_in_activate),
    .io_in_weight(PE_Array_4_7_io_in_weight),
    .io_in_psum(PE_Array_4_7_io_in_psum),
    .io_in_flow(PE_Array_4_7_io_in_flow),
    .io_in_shift(PE_Array_4_7_io_in_shift),
    .io_out_activate(PE_Array_4_7_io_out_activate),
    .io_out_weight(PE_Array_4_7_io_out_weight),
    .io_out_psum(PE_Array_4_7_io_out_psum)
  );
  basic_PE PE_Array_4_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_8_clock),
    .reset(PE_Array_4_8_reset),
    .io_in_activate(PE_Array_4_8_io_in_activate),
    .io_in_weight(PE_Array_4_8_io_in_weight),
    .io_in_psum(PE_Array_4_8_io_in_psum),
    .io_in_flow(PE_Array_4_8_io_in_flow),
    .io_in_shift(PE_Array_4_8_io_in_shift),
    .io_out_activate(PE_Array_4_8_io_out_activate),
    .io_out_weight(PE_Array_4_8_io_out_weight),
    .io_out_psum(PE_Array_4_8_io_out_psum)
  );
  basic_PE PE_Array_4_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_9_clock),
    .reset(PE_Array_4_9_reset),
    .io_in_activate(PE_Array_4_9_io_in_activate),
    .io_in_weight(PE_Array_4_9_io_in_weight),
    .io_in_psum(PE_Array_4_9_io_in_psum),
    .io_in_flow(PE_Array_4_9_io_in_flow),
    .io_in_shift(PE_Array_4_9_io_in_shift),
    .io_out_activate(PE_Array_4_9_io_out_activate),
    .io_out_weight(PE_Array_4_9_io_out_weight),
    .io_out_psum(PE_Array_4_9_io_out_psum)
  );
  basic_PE PE_Array_4_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_10_clock),
    .reset(PE_Array_4_10_reset),
    .io_in_activate(PE_Array_4_10_io_in_activate),
    .io_in_weight(PE_Array_4_10_io_in_weight),
    .io_in_psum(PE_Array_4_10_io_in_psum),
    .io_in_flow(PE_Array_4_10_io_in_flow),
    .io_in_shift(PE_Array_4_10_io_in_shift),
    .io_out_activate(PE_Array_4_10_io_out_activate),
    .io_out_weight(PE_Array_4_10_io_out_weight),
    .io_out_psum(PE_Array_4_10_io_out_psum)
  );
  basic_PE PE_Array_4_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_11_clock),
    .reset(PE_Array_4_11_reset),
    .io_in_activate(PE_Array_4_11_io_in_activate),
    .io_in_weight(PE_Array_4_11_io_in_weight),
    .io_in_psum(PE_Array_4_11_io_in_psum),
    .io_in_flow(PE_Array_4_11_io_in_flow),
    .io_in_shift(PE_Array_4_11_io_in_shift),
    .io_out_activate(PE_Array_4_11_io_out_activate),
    .io_out_weight(PE_Array_4_11_io_out_weight),
    .io_out_psum(PE_Array_4_11_io_out_psum)
  );
  basic_PE PE_Array_4_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_12_clock),
    .reset(PE_Array_4_12_reset),
    .io_in_activate(PE_Array_4_12_io_in_activate),
    .io_in_weight(PE_Array_4_12_io_in_weight),
    .io_in_psum(PE_Array_4_12_io_in_psum),
    .io_in_flow(PE_Array_4_12_io_in_flow),
    .io_in_shift(PE_Array_4_12_io_in_shift),
    .io_out_activate(PE_Array_4_12_io_out_activate),
    .io_out_weight(PE_Array_4_12_io_out_weight),
    .io_out_psum(PE_Array_4_12_io_out_psum)
  );
  basic_PE PE_Array_4_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_13_clock),
    .reset(PE_Array_4_13_reset),
    .io_in_activate(PE_Array_4_13_io_in_activate),
    .io_in_weight(PE_Array_4_13_io_in_weight),
    .io_in_psum(PE_Array_4_13_io_in_psum),
    .io_in_flow(PE_Array_4_13_io_in_flow),
    .io_in_shift(PE_Array_4_13_io_in_shift),
    .io_out_activate(PE_Array_4_13_io_out_activate),
    .io_out_weight(PE_Array_4_13_io_out_weight),
    .io_out_psum(PE_Array_4_13_io_out_psum)
  );
  basic_PE PE_Array_4_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_14_clock),
    .reset(PE_Array_4_14_reset),
    .io_in_activate(PE_Array_4_14_io_in_activate),
    .io_in_weight(PE_Array_4_14_io_in_weight),
    .io_in_psum(PE_Array_4_14_io_in_psum),
    .io_in_flow(PE_Array_4_14_io_in_flow),
    .io_in_shift(PE_Array_4_14_io_in_shift),
    .io_out_activate(PE_Array_4_14_io_out_activate),
    .io_out_weight(PE_Array_4_14_io_out_weight),
    .io_out_psum(PE_Array_4_14_io_out_psum)
  );
  basic_PE PE_Array_4_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_15_clock),
    .reset(PE_Array_4_15_reset),
    .io_in_activate(PE_Array_4_15_io_in_activate),
    .io_in_weight(PE_Array_4_15_io_in_weight),
    .io_in_psum(PE_Array_4_15_io_in_psum),
    .io_in_flow(PE_Array_4_15_io_in_flow),
    .io_in_shift(PE_Array_4_15_io_in_shift),
    .io_out_activate(PE_Array_4_15_io_out_activate),
    .io_out_weight(PE_Array_4_15_io_out_weight),
    .io_out_psum(PE_Array_4_15_io_out_psum)
  );
  basic_PE PE_Array_5_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_0_clock),
    .reset(PE_Array_5_0_reset),
    .io_in_activate(PE_Array_5_0_io_in_activate),
    .io_in_weight(PE_Array_5_0_io_in_weight),
    .io_in_psum(PE_Array_5_0_io_in_psum),
    .io_in_flow(PE_Array_5_0_io_in_flow),
    .io_in_shift(PE_Array_5_0_io_in_shift),
    .io_out_activate(PE_Array_5_0_io_out_activate),
    .io_out_weight(PE_Array_5_0_io_out_weight),
    .io_out_psum(PE_Array_5_0_io_out_psum)
  );
  basic_PE PE_Array_5_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_1_clock),
    .reset(PE_Array_5_1_reset),
    .io_in_activate(PE_Array_5_1_io_in_activate),
    .io_in_weight(PE_Array_5_1_io_in_weight),
    .io_in_psum(PE_Array_5_1_io_in_psum),
    .io_in_flow(PE_Array_5_1_io_in_flow),
    .io_in_shift(PE_Array_5_1_io_in_shift),
    .io_out_activate(PE_Array_5_1_io_out_activate),
    .io_out_weight(PE_Array_5_1_io_out_weight),
    .io_out_psum(PE_Array_5_1_io_out_psum)
  );
  basic_PE PE_Array_5_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_2_clock),
    .reset(PE_Array_5_2_reset),
    .io_in_activate(PE_Array_5_2_io_in_activate),
    .io_in_weight(PE_Array_5_2_io_in_weight),
    .io_in_psum(PE_Array_5_2_io_in_psum),
    .io_in_flow(PE_Array_5_2_io_in_flow),
    .io_in_shift(PE_Array_5_2_io_in_shift),
    .io_out_activate(PE_Array_5_2_io_out_activate),
    .io_out_weight(PE_Array_5_2_io_out_weight),
    .io_out_psum(PE_Array_5_2_io_out_psum)
  );
  basic_PE PE_Array_5_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_3_clock),
    .reset(PE_Array_5_3_reset),
    .io_in_activate(PE_Array_5_3_io_in_activate),
    .io_in_weight(PE_Array_5_3_io_in_weight),
    .io_in_psum(PE_Array_5_3_io_in_psum),
    .io_in_flow(PE_Array_5_3_io_in_flow),
    .io_in_shift(PE_Array_5_3_io_in_shift),
    .io_out_activate(PE_Array_5_3_io_out_activate),
    .io_out_weight(PE_Array_5_3_io_out_weight),
    .io_out_psum(PE_Array_5_3_io_out_psum)
  );
  basic_PE PE_Array_5_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_4_clock),
    .reset(PE_Array_5_4_reset),
    .io_in_activate(PE_Array_5_4_io_in_activate),
    .io_in_weight(PE_Array_5_4_io_in_weight),
    .io_in_psum(PE_Array_5_4_io_in_psum),
    .io_in_flow(PE_Array_5_4_io_in_flow),
    .io_in_shift(PE_Array_5_4_io_in_shift),
    .io_out_activate(PE_Array_5_4_io_out_activate),
    .io_out_weight(PE_Array_5_4_io_out_weight),
    .io_out_psum(PE_Array_5_4_io_out_psum)
  );
  basic_PE PE_Array_5_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_5_clock),
    .reset(PE_Array_5_5_reset),
    .io_in_activate(PE_Array_5_5_io_in_activate),
    .io_in_weight(PE_Array_5_5_io_in_weight),
    .io_in_psum(PE_Array_5_5_io_in_psum),
    .io_in_flow(PE_Array_5_5_io_in_flow),
    .io_in_shift(PE_Array_5_5_io_in_shift),
    .io_out_activate(PE_Array_5_5_io_out_activate),
    .io_out_weight(PE_Array_5_5_io_out_weight),
    .io_out_psum(PE_Array_5_5_io_out_psum)
  );
  basic_PE PE_Array_5_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_6_clock),
    .reset(PE_Array_5_6_reset),
    .io_in_activate(PE_Array_5_6_io_in_activate),
    .io_in_weight(PE_Array_5_6_io_in_weight),
    .io_in_psum(PE_Array_5_6_io_in_psum),
    .io_in_flow(PE_Array_5_6_io_in_flow),
    .io_in_shift(PE_Array_5_6_io_in_shift),
    .io_out_activate(PE_Array_5_6_io_out_activate),
    .io_out_weight(PE_Array_5_6_io_out_weight),
    .io_out_psum(PE_Array_5_6_io_out_psum)
  );
  basic_PE PE_Array_5_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_7_clock),
    .reset(PE_Array_5_7_reset),
    .io_in_activate(PE_Array_5_7_io_in_activate),
    .io_in_weight(PE_Array_5_7_io_in_weight),
    .io_in_psum(PE_Array_5_7_io_in_psum),
    .io_in_flow(PE_Array_5_7_io_in_flow),
    .io_in_shift(PE_Array_5_7_io_in_shift),
    .io_out_activate(PE_Array_5_7_io_out_activate),
    .io_out_weight(PE_Array_5_7_io_out_weight),
    .io_out_psum(PE_Array_5_7_io_out_psum)
  );
  basic_PE PE_Array_5_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_8_clock),
    .reset(PE_Array_5_8_reset),
    .io_in_activate(PE_Array_5_8_io_in_activate),
    .io_in_weight(PE_Array_5_8_io_in_weight),
    .io_in_psum(PE_Array_5_8_io_in_psum),
    .io_in_flow(PE_Array_5_8_io_in_flow),
    .io_in_shift(PE_Array_5_8_io_in_shift),
    .io_out_activate(PE_Array_5_8_io_out_activate),
    .io_out_weight(PE_Array_5_8_io_out_weight),
    .io_out_psum(PE_Array_5_8_io_out_psum)
  );
  basic_PE PE_Array_5_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_9_clock),
    .reset(PE_Array_5_9_reset),
    .io_in_activate(PE_Array_5_9_io_in_activate),
    .io_in_weight(PE_Array_5_9_io_in_weight),
    .io_in_psum(PE_Array_5_9_io_in_psum),
    .io_in_flow(PE_Array_5_9_io_in_flow),
    .io_in_shift(PE_Array_5_9_io_in_shift),
    .io_out_activate(PE_Array_5_9_io_out_activate),
    .io_out_weight(PE_Array_5_9_io_out_weight),
    .io_out_psum(PE_Array_5_9_io_out_psum)
  );
  basic_PE PE_Array_5_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_10_clock),
    .reset(PE_Array_5_10_reset),
    .io_in_activate(PE_Array_5_10_io_in_activate),
    .io_in_weight(PE_Array_5_10_io_in_weight),
    .io_in_psum(PE_Array_5_10_io_in_psum),
    .io_in_flow(PE_Array_5_10_io_in_flow),
    .io_in_shift(PE_Array_5_10_io_in_shift),
    .io_out_activate(PE_Array_5_10_io_out_activate),
    .io_out_weight(PE_Array_5_10_io_out_weight),
    .io_out_psum(PE_Array_5_10_io_out_psum)
  );
  basic_PE PE_Array_5_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_11_clock),
    .reset(PE_Array_5_11_reset),
    .io_in_activate(PE_Array_5_11_io_in_activate),
    .io_in_weight(PE_Array_5_11_io_in_weight),
    .io_in_psum(PE_Array_5_11_io_in_psum),
    .io_in_flow(PE_Array_5_11_io_in_flow),
    .io_in_shift(PE_Array_5_11_io_in_shift),
    .io_out_activate(PE_Array_5_11_io_out_activate),
    .io_out_weight(PE_Array_5_11_io_out_weight),
    .io_out_psum(PE_Array_5_11_io_out_psum)
  );
  basic_PE PE_Array_5_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_12_clock),
    .reset(PE_Array_5_12_reset),
    .io_in_activate(PE_Array_5_12_io_in_activate),
    .io_in_weight(PE_Array_5_12_io_in_weight),
    .io_in_psum(PE_Array_5_12_io_in_psum),
    .io_in_flow(PE_Array_5_12_io_in_flow),
    .io_in_shift(PE_Array_5_12_io_in_shift),
    .io_out_activate(PE_Array_5_12_io_out_activate),
    .io_out_weight(PE_Array_5_12_io_out_weight),
    .io_out_psum(PE_Array_5_12_io_out_psum)
  );
  basic_PE PE_Array_5_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_13_clock),
    .reset(PE_Array_5_13_reset),
    .io_in_activate(PE_Array_5_13_io_in_activate),
    .io_in_weight(PE_Array_5_13_io_in_weight),
    .io_in_psum(PE_Array_5_13_io_in_psum),
    .io_in_flow(PE_Array_5_13_io_in_flow),
    .io_in_shift(PE_Array_5_13_io_in_shift),
    .io_out_activate(PE_Array_5_13_io_out_activate),
    .io_out_weight(PE_Array_5_13_io_out_weight),
    .io_out_psum(PE_Array_5_13_io_out_psum)
  );
  basic_PE PE_Array_5_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_14_clock),
    .reset(PE_Array_5_14_reset),
    .io_in_activate(PE_Array_5_14_io_in_activate),
    .io_in_weight(PE_Array_5_14_io_in_weight),
    .io_in_psum(PE_Array_5_14_io_in_psum),
    .io_in_flow(PE_Array_5_14_io_in_flow),
    .io_in_shift(PE_Array_5_14_io_in_shift),
    .io_out_activate(PE_Array_5_14_io_out_activate),
    .io_out_weight(PE_Array_5_14_io_out_weight),
    .io_out_psum(PE_Array_5_14_io_out_psum)
  );
  basic_PE PE_Array_5_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_15_clock),
    .reset(PE_Array_5_15_reset),
    .io_in_activate(PE_Array_5_15_io_in_activate),
    .io_in_weight(PE_Array_5_15_io_in_weight),
    .io_in_psum(PE_Array_5_15_io_in_psum),
    .io_in_flow(PE_Array_5_15_io_in_flow),
    .io_in_shift(PE_Array_5_15_io_in_shift),
    .io_out_activate(PE_Array_5_15_io_out_activate),
    .io_out_weight(PE_Array_5_15_io_out_weight),
    .io_out_psum(PE_Array_5_15_io_out_psum)
  );
  basic_PE PE_Array_6_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_0_clock),
    .reset(PE_Array_6_0_reset),
    .io_in_activate(PE_Array_6_0_io_in_activate),
    .io_in_weight(PE_Array_6_0_io_in_weight),
    .io_in_psum(PE_Array_6_0_io_in_psum),
    .io_in_flow(PE_Array_6_0_io_in_flow),
    .io_in_shift(PE_Array_6_0_io_in_shift),
    .io_out_activate(PE_Array_6_0_io_out_activate),
    .io_out_weight(PE_Array_6_0_io_out_weight),
    .io_out_psum(PE_Array_6_0_io_out_psum)
  );
  basic_PE PE_Array_6_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_1_clock),
    .reset(PE_Array_6_1_reset),
    .io_in_activate(PE_Array_6_1_io_in_activate),
    .io_in_weight(PE_Array_6_1_io_in_weight),
    .io_in_psum(PE_Array_6_1_io_in_psum),
    .io_in_flow(PE_Array_6_1_io_in_flow),
    .io_in_shift(PE_Array_6_1_io_in_shift),
    .io_out_activate(PE_Array_6_1_io_out_activate),
    .io_out_weight(PE_Array_6_1_io_out_weight),
    .io_out_psum(PE_Array_6_1_io_out_psum)
  );
  basic_PE PE_Array_6_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_2_clock),
    .reset(PE_Array_6_2_reset),
    .io_in_activate(PE_Array_6_2_io_in_activate),
    .io_in_weight(PE_Array_6_2_io_in_weight),
    .io_in_psum(PE_Array_6_2_io_in_psum),
    .io_in_flow(PE_Array_6_2_io_in_flow),
    .io_in_shift(PE_Array_6_2_io_in_shift),
    .io_out_activate(PE_Array_6_2_io_out_activate),
    .io_out_weight(PE_Array_6_2_io_out_weight),
    .io_out_psum(PE_Array_6_2_io_out_psum)
  );
  basic_PE PE_Array_6_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_3_clock),
    .reset(PE_Array_6_3_reset),
    .io_in_activate(PE_Array_6_3_io_in_activate),
    .io_in_weight(PE_Array_6_3_io_in_weight),
    .io_in_psum(PE_Array_6_3_io_in_psum),
    .io_in_flow(PE_Array_6_3_io_in_flow),
    .io_in_shift(PE_Array_6_3_io_in_shift),
    .io_out_activate(PE_Array_6_3_io_out_activate),
    .io_out_weight(PE_Array_6_3_io_out_weight),
    .io_out_psum(PE_Array_6_3_io_out_psum)
  );
  basic_PE PE_Array_6_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_4_clock),
    .reset(PE_Array_6_4_reset),
    .io_in_activate(PE_Array_6_4_io_in_activate),
    .io_in_weight(PE_Array_6_4_io_in_weight),
    .io_in_psum(PE_Array_6_4_io_in_psum),
    .io_in_flow(PE_Array_6_4_io_in_flow),
    .io_in_shift(PE_Array_6_4_io_in_shift),
    .io_out_activate(PE_Array_6_4_io_out_activate),
    .io_out_weight(PE_Array_6_4_io_out_weight),
    .io_out_psum(PE_Array_6_4_io_out_psum)
  );
  basic_PE PE_Array_6_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_5_clock),
    .reset(PE_Array_6_5_reset),
    .io_in_activate(PE_Array_6_5_io_in_activate),
    .io_in_weight(PE_Array_6_5_io_in_weight),
    .io_in_psum(PE_Array_6_5_io_in_psum),
    .io_in_flow(PE_Array_6_5_io_in_flow),
    .io_in_shift(PE_Array_6_5_io_in_shift),
    .io_out_activate(PE_Array_6_5_io_out_activate),
    .io_out_weight(PE_Array_6_5_io_out_weight),
    .io_out_psum(PE_Array_6_5_io_out_psum)
  );
  basic_PE PE_Array_6_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_6_clock),
    .reset(PE_Array_6_6_reset),
    .io_in_activate(PE_Array_6_6_io_in_activate),
    .io_in_weight(PE_Array_6_6_io_in_weight),
    .io_in_psum(PE_Array_6_6_io_in_psum),
    .io_in_flow(PE_Array_6_6_io_in_flow),
    .io_in_shift(PE_Array_6_6_io_in_shift),
    .io_out_activate(PE_Array_6_6_io_out_activate),
    .io_out_weight(PE_Array_6_6_io_out_weight),
    .io_out_psum(PE_Array_6_6_io_out_psum)
  );
  basic_PE PE_Array_6_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_7_clock),
    .reset(PE_Array_6_7_reset),
    .io_in_activate(PE_Array_6_7_io_in_activate),
    .io_in_weight(PE_Array_6_7_io_in_weight),
    .io_in_psum(PE_Array_6_7_io_in_psum),
    .io_in_flow(PE_Array_6_7_io_in_flow),
    .io_in_shift(PE_Array_6_7_io_in_shift),
    .io_out_activate(PE_Array_6_7_io_out_activate),
    .io_out_weight(PE_Array_6_7_io_out_weight),
    .io_out_psum(PE_Array_6_7_io_out_psum)
  );
  basic_PE PE_Array_6_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_8_clock),
    .reset(PE_Array_6_8_reset),
    .io_in_activate(PE_Array_6_8_io_in_activate),
    .io_in_weight(PE_Array_6_8_io_in_weight),
    .io_in_psum(PE_Array_6_8_io_in_psum),
    .io_in_flow(PE_Array_6_8_io_in_flow),
    .io_in_shift(PE_Array_6_8_io_in_shift),
    .io_out_activate(PE_Array_6_8_io_out_activate),
    .io_out_weight(PE_Array_6_8_io_out_weight),
    .io_out_psum(PE_Array_6_8_io_out_psum)
  );
  basic_PE PE_Array_6_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_9_clock),
    .reset(PE_Array_6_9_reset),
    .io_in_activate(PE_Array_6_9_io_in_activate),
    .io_in_weight(PE_Array_6_9_io_in_weight),
    .io_in_psum(PE_Array_6_9_io_in_psum),
    .io_in_flow(PE_Array_6_9_io_in_flow),
    .io_in_shift(PE_Array_6_9_io_in_shift),
    .io_out_activate(PE_Array_6_9_io_out_activate),
    .io_out_weight(PE_Array_6_9_io_out_weight),
    .io_out_psum(PE_Array_6_9_io_out_psum)
  );
  basic_PE PE_Array_6_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_10_clock),
    .reset(PE_Array_6_10_reset),
    .io_in_activate(PE_Array_6_10_io_in_activate),
    .io_in_weight(PE_Array_6_10_io_in_weight),
    .io_in_psum(PE_Array_6_10_io_in_psum),
    .io_in_flow(PE_Array_6_10_io_in_flow),
    .io_in_shift(PE_Array_6_10_io_in_shift),
    .io_out_activate(PE_Array_6_10_io_out_activate),
    .io_out_weight(PE_Array_6_10_io_out_weight),
    .io_out_psum(PE_Array_6_10_io_out_psum)
  );
  basic_PE PE_Array_6_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_11_clock),
    .reset(PE_Array_6_11_reset),
    .io_in_activate(PE_Array_6_11_io_in_activate),
    .io_in_weight(PE_Array_6_11_io_in_weight),
    .io_in_psum(PE_Array_6_11_io_in_psum),
    .io_in_flow(PE_Array_6_11_io_in_flow),
    .io_in_shift(PE_Array_6_11_io_in_shift),
    .io_out_activate(PE_Array_6_11_io_out_activate),
    .io_out_weight(PE_Array_6_11_io_out_weight),
    .io_out_psum(PE_Array_6_11_io_out_psum)
  );
  basic_PE PE_Array_6_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_12_clock),
    .reset(PE_Array_6_12_reset),
    .io_in_activate(PE_Array_6_12_io_in_activate),
    .io_in_weight(PE_Array_6_12_io_in_weight),
    .io_in_psum(PE_Array_6_12_io_in_psum),
    .io_in_flow(PE_Array_6_12_io_in_flow),
    .io_in_shift(PE_Array_6_12_io_in_shift),
    .io_out_activate(PE_Array_6_12_io_out_activate),
    .io_out_weight(PE_Array_6_12_io_out_weight),
    .io_out_psum(PE_Array_6_12_io_out_psum)
  );
  basic_PE PE_Array_6_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_13_clock),
    .reset(PE_Array_6_13_reset),
    .io_in_activate(PE_Array_6_13_io_in_activate),
    .io_in_weight(PE_Array_6_13_io_in_weight),
    .io_in_psum(PE_Array_6_13_io_in_psum),
    .io_in_flow(PE_Array_6_13_io_in_flow),
    .io_in_shift(PE_Array_6_13_io_in_shift),
    .io_out_activate(PE_Array_6_13_io_out_activate),
    .io_out_weight(PE_Array_6_13_io_out_weight),
    .io_out_psum(PE_Array_6_13_io_out_psum)
  );
  basic_PE PE_Array_6_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_14_clock),
    .reset(PE_Array_6_14_reset),
    .io_in_activate(PE_Array_6_14_io_in_activate),
    .io_in_weight(PE_Array_6_14_io_in_weight),
    .io_in_psum(PE_Array_6_14_io_in_psum),
    .io_in_flow(PE_Array_6_14_io_in_flow),
    .io_in_shift(PE_Array_6_14_io_in_shift),
    .io_out_activate(PE_Array_6_14_io_out_activate),
    .io_out_weight(PE_Array_6_14_io_out_weight),
    .io_out_psum(PE_Array_6_14_io_out_psum)
  );
  basic_PE PE_Array_6_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_15_clock),
    .reset(PE_Array_6_15_reset),
    .io_in_activate(PE_Array_6_15_io_in_activate),
    .io_in_weight(PE_Array_6_15_io_in_weight),
    .io_in_psum(PE_Array_6_15_io_in_psum),
    .io_in_flow(PE_Array_6_15_io_in_flow),
    .io_in_shift(PE_Array_6_15_io_in_shift),
    .io_out_activate(PE_Array_6_15_io_out_activate),
    .io_out_weight(PE_Array_6_15_io_out_weight),
    .io_out_psum(PE_Array_6_15_io_out_psum)
  );
  basic_PE PE_Array_7_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_0_clock),
    .reset(PE_Array_7_0_reset),
    .io_in_activate(PE_Array_7_0_io_in_activate),
    .io_in_weight(PE_Array_7_0_io_in_weight),
    .io_in_psum(PE_Array_7_0_io_in_psum),
    .io_in_flow(PE_Array_7_0_io_in_flow),
    .io_in_shift(PE_Array_7_0_io_in_shift),
    .io_out_activate(PE_Array_7_0_io_out_activate),
    .io_out_weight(PE_Array_7_0_io_out_weight),
    .io_out_psum(PE_Array_7_0_io_out_psum)
  );
  basic_PE PE_Array_7_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_1_clock),
    .reset(PE_Array_7_1_reset),
    .io_in_activate(PE_Array_7_1_io_in_activate),
    .io_in_weight(PE_Array_7_1_io_in_weight),
    .io_in_psum(PE_Array_7_1_io_in_psum),
    .io_in_flow(PE_Array_7_1_io_in_flow),
    .io_in_shift(PE_Array_7_1_io_in_shift),
    .io_out_activate(PE_Array_7_1_io_out_activate),
    .io_out_weight(PE_Array_7_1_io_out_weight),
    .io_out_psum(PE_Array_7_1_io_out_psum)
  );
  basic_PE PE_Array_7_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_2_clock),
    .reset(PE_Array_7_2_reset),
    .io_in_activate(PE_Array_7_2_io_in_activate),
    .io_in_weight(PE_Array_7_2_io_in_weight),
    .io_in_psum(PE_Array_7_2_io_in_psum),
    .io_in_flow(PE_Array_7_2_io_in_flow),
    .io_in_shift(PE_Array_7_2_io_in_shift),
    .io_out_activate(PE_Array_7_2_io_out_activate),
    .io_out_weight(PE_Array_7_2_io_out_weight),
    .io_out_psum(PE_Array_7_2_io_out_psum)
  );
  basic_PE PE_Array_7_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_3_clock),
    .reset(PE_Array_7_3_reset),
    .io_in_activate(PE_Array_7_3_io_in_activate),
    .io_in_weight(PE_Array_7_3_io_in_weight),
    .io_in_psum(PE_Array_7_3_io_in_psum),
    .io_in_flow(PE_Array_7_3_io_in_flow),
    .io_in_shift(PE_Array_7_3_io_in_shift),
    .io_out_activate(PE_Array_7_3_io_out_activate),
    .io_out_weight(PE_Array_7_3_io_out_weight),
    .io_out_psum(PE_Array_7_3_io_out_psum)
  );
  basic_PE PE_Array_7_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_4_clock),
    .reset(PE_Array_7_4_reset),
    .io_in_activate(PE_Array_7_4_io_in_activate),
    .io_in_weight(PE_Array_7_4_io_in_weight),
    .io_in_psum(PE_Array_7_4_io_in_psum),
    .io_in_flow(PE_Array_7_4_io_in_flow),
    .io_in_shift(PE_Array_7_4_io_in_shift),
    .io_out_activate(PE_Array_7_4_io_out_activate),
    .io_out_weight(PE_Array_7_4_io_out_weight),
    .io_out_psum(PE_Array_7_4_io_out_psum)
  );
  basic_PE PE_Array_7_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_5_clock),
    .reset(PE_Array_7_5_reset),
    .io_in_activate(PE_Array_7_5_io_in_activate),
    .io_in_weight(PE_Array_7_5_io_in_weight),
    .io_in_psum(PE_Array_7_5_io_in_psum),
    .io_in_flow(PE_Array_7_5_io_in_flow),
    .io_in_shift(PE_Array_7_5_io_in_shift),
    .io_out_activate(PE_Array_7_5_io_out_activate),
    .io_out_weight(PE_Array_7_5_io_out_weight),
    .io_out_psum(PE_Array_7_5_io_out_psum)
  );
  basic_PE PE_Array_7_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_6_clock),
    .reset(PE_Array_7_6_reset),
    .io_in_activate(PE_Array_7_6_io_in_activate),
    .io_in_weight(PE_Array_7_6_io_in_weight),
    .io_in_psum(PE_Array_7_6_io_in_psum),
    .io_in_flow(PE_Array_7_6_io_in_flow),
    .io_in_shift(PE_Array_7_6_io_in_shift),
    .io_out_activate(PE_Array_7_6_io_out_activate),
    .io_out_weight(PE_Array_7_6_io_out_weight),
    .io_out_psum(PE_Array_7_6_io_out_psum)
  );
  basic_PE PE_Array_7_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_7_clock),
    .reset(PE_Array_7_7_reset),
    .io_in_activate(PE_Array_7_7_io_in_activate),
    .io_in_weight(PE_Array_7_7_io_in_weight),
    .io_in_psum(PE_Array_7_7_io_in_psum),
    .io_in_flow(PE_Array_7_7_io_in_flow),
    .io_in_shift(PE_Array_7_7_io_in_shift),
    .io_out_activate(PE_Array_7_7_io_out_activate),
    .io_out_weight(PE_Array_7_7_io_out_weight),
    .io_out_psum(PE_Array_7_7_io_out_psum)
  );
  basic_PE PE_Array_7_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_8_clock),
    .reset(PE_Array_7_8_reset),
    .io_in_activate(PE_Array_7_8_io_in_activate),
    .io_in_weight(PE_Array_7_8_io_in_weight),
    .io_in_psum(PE_Array_7_8_io_in_psum),
    .io_in_flow(PE_Array_7_8_io_in_flow),
    .io_in_shift(PE_Array_7_8_io_in_shift),
    .io_out_activate(PE_Array_7_8_io_out_activate),
    .io_out_weight(PE_Array_7_8_io_out_weight),
    .io_out_psum(PE_Array_7_8_io_out_psum)
  );
  basic_PE PE_Array_7_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_9_clock),
    .reset(PE_Array_7_9_reset),
    .io_in_activate(PE_Array_7_9_io_in_activate),
    .io_in_weight(PE_Array_7_9_io_in_weight),
    .io_in_psum(PE_Array_7_9_io_in_psum),
    .io_in_flow(PE_Array_7_9_io_in_flow),
    .io_in_shift(PE_Array_7_9_io_in_shift),
    .io_out_activate(PE_Array_7_9_io_out_activate),
    .io_out_weight(PE_Array_7_9_io_out_weight),
    .io_out_psum(PE_Array_7_9_io_out_psum)
  );
  basic_PE PE_Array_7_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_10_clock),
    .reset(PE_Array_7_10_reset),
    .io_in_activate(PE_Array_7_10_io_in_activate),
    .io_in_weight(PE_Array_7_10_io_in_weight),
    .io_in_psum(PE_Array_7_10_io_in_psum),
    .io_in_flow(PE_Array_7_10_io_in_flow),
    .io_in_shift(PE_Array_7_10_io_in_shift),
    .io_out_activate(PE_Array_7_10_io_out_activate),
    .io_out_weight(PE_Array_7_10_io_out_weight),
    .io_out_psum(PE_Array_7_10_io_out_psum)
  );
  basic_PE PE_Array_7_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_11_clock),
    .reset(PE_Array_7_11_reset),
    .io_in_activate(PE_Array_7_11_io_in_activate),
    .io_in_weight(PE_Array_7_11_io_in_weight),
    .io_in_psum(PE_Array_7_11_io_in_psum),
    .io_in_flow(PE_Array_7_11_io_in_flow),
    .io_in_shift(PE_Array_7_11_io_in_shift),
    .io_out_activate(PE_Array_7_11_io_out_activate),
    .io_out_weight(PE_Array_7_11_io_out_weight),
    .io_out_psum(PE_Array_7_11_io_out_psum)
  );
  basic_PE PE_Array_7_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_12_clock),
    .reset(PE_Array_7_12_reset),
    .io_in_activate(PE_Array_7_12_io_in_activate),
    .io_in_weight(PE_Array_7_12_io_in_weight),
    .io_in_psum(PE_Array_7_12_io_in_psum),
    .io_in_flow(PE_Array_7_12_io_in_flow),
    .io_in_shift(PE_Array_7_12_io_in_shift),
    .io_out_activate(PE_Array_7_12_io_out_activate),
    .io_out_weight(PE_Array_7_12_io_out_weight),
    .io_out_psum(PE_Array_7_12_io_out_psum)
  );
  basic_PE PE_Array_7_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_13_clock),
    .reset(PE_Array_7_13_reset),
    .io_in_activate(PE_Array_7_13_io_in_activate),
    .io_in_weight(PE_Array_7_13_io_in_weight),
    .io_in_psum(PE_Array_7_13_io_in_psum),
    .io_in_flow(PE_Array_7_13_io_in_flow),
    .io_in_shift(PE_Array_7_13_io_in_shift),
    .io_out_activate(PE_Array_7_13_io_out_activate),
    .io_out_weight(PE_Array_7_13_io_out_weight),
    .io_out_psum(PE_Array_7_13_io_out_psum)
  );
  basic_PE PE_Array_7_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_14_clock),
    .reset(PE_Array_7_14_reset),
    .io_in_activate(PE_Array_7_14_io_in_activate),
    .io_in_weight(PE_Array_7_14_io_in_weight),
    .io_in_psum(PE_Array_7_14_io_in_psum),
    .io_in_flow(PE_Array_7_14_io_in_flow),
    .io_in_shift(PE_Array_7_14_io_in_shift),
    .io_out_activate(PE_Array_7_14_io_out_activate),
    .io_out_weight(PE_Array_7_14_io_out_weight),
    .io_out_psum(PE_Array_7_14_io_out_psum)
  );
  basic_PE PE_Array_7_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_15_clock),
    .reset(PE_Array_7_15_reset),
    .io_in_activate(PE_Array_7_15_io_in_activate),
    .io_in_weight(PE_Array_7_15_io_in_weight),
    .io_in_psum(PE_Array_7_15_io_in_psum),
    .io_in_flow(PE_Array_7_15_io_in_flow),
    .io_in_shift(PE_Array_7_15_io_in_shift),
    .io_out_activate(PE_Array_7_15_io_out_activate),
    .io_out_weight(PE_Array_7_15_io_out_weight),
    .io_out_psum(PE_Array_7_15_io_out_psum)
  );
  basic_PE PE_Array_8_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_0_clock),
    .reset(PE_Array_8_0_reset),
    .io_in_activate(PE_Array_8_0_io_in_activate),
    .io_in_weight(PE_Array_8_0_io_in_weight),
    .io_in_psum(PE_Array_8_0_io_in_psum),
    .io_in_flow(PE_Array_8_0_io_in_flow),
    .io_in_shift(PE_Array_8_0_io_in_shift),
    .io_out_activate(PE_Array_8_0_io_out_activate),
    .io_out_weight(PE_Array_8_0_io_out_weight),
    .io_out_psum(PE_Array_8_0_io_out_psum)
  );
  basic_PE PE_Array_8_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_1_clock),
    .reset(PE_Array_8_1_reset),
    .io_in_activate(PE_Array_8_1_io_in_activate),
    .io_in_weight(PE_Array_8_1_io_in_weight),
    .io_in_psum(PE_Array_8_1_io_in_psum),
    .io_in_flow(PE_Array_8_1_io_in_flow),
    .io_in_shift(PE_Array_8_1_io_in_shift),
    .io_out_activate(PE_Array_8_1_io_out_activate),
    .io_out_weight(PE_Array_8_1_io_out_weight),
    .io_out_psum(PE_Array_8_1_io_out_psum)
  );
  basic_PE PE_Array_8_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_2_clock),
    .reset(PE_Array_8_2_reset),
    .io_in_activate(PE_Array_8_2_io_in_activate),
    .io_in_weight(PE_Array_8_2_io_in_weight),
    .io_in_psum(PE_Array_8_2_io_in_psum),
    .io_in_flow(PE_Array_8_2_io_in_flow),
    .io_in_shift(PE_Array_8_2_io_in_shift),
    .io_out_activate(PE_Array_8_2_io_out_activate),
    .io_out_weight(PE_Array_8_2_io_out_weight),
    .io_out_psum(PE_Array_8_2_io_out_psum)
  );
  basic_PE PE_Array_8_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_3_clock),
    .reset(PE_Array_8_3_reset),
    .io_in_activate(PE_Array_8_3_io_in_activate),
    .io_in_weight(PE_Array_8_3_io_in_weight),
    .io_in_psum(PE_Array_8_3_io_in_psum),
    .io_in_flow(PE_Array_8_3_io_in_flow),
    .io_in_shift(PE_Array_8_3_io_in_shift),
    .io_out_activate(PE_Array_8_3_io_out_activate),
    .io_out_weight(PE_Array_8_3_io_out_weight),
    .io_out_psum(PE_Array_8_3_io_out_psum)
  );
  basic_PE PE_Array_8_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_4_clock),
    .reset(PE_Array_8_4_reset),
    .io_in_activate(PE_Array_8_4_io_in_activate),
    .io_in_weight(PE_Array_8_4_io_in_weight),
    .io_in_psum(PE_Array_8_4_io_in_psum),
    .io_in_flow(PE_Array_8_4_io_in_flow),
    .io_in_shift(PE_Array_8_4_io_in_shift),
    .io_out_activate(PE_Array_8_4_io_out_activate),
    .io_out_weight(PE_Array_8_4_io_out_weight),
    .io_out_psum(PE_Array_8_4_io_out_psum)
  );
  basic_PE PE_Array_8_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_5_clock),
    .reset(PE_Array_8_5_reset),
    .io_in_activate(PE_Array_8_5_io_in_activate),
    .io_in_weight(PE_Array_8_5_io_in_weight),
    .io_in_psum(PE_Array_8_5_io_in_psum),
    .io_in_flow(PE_Array_8_5_io_in_flow),
    .io_in_shift(PE_Array_8_5_io_in_shift),
    .io_out_activate(PE_Array_8_5_io_out_activate),
    .io_out_weight(PE_Array_8_5_io_out_weight),
    .io_out_psum(PE_Array_8_5_io_out_psum)
  );
  basic_PE PE_Array_8_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_6_clock),
    .reset(PE_Array_8_6_reset),
    .io_in_activate(PE_Array_8_6_io_in_activate),
    .io_in_weight(PE_Array_8_6_io_in_weight),
    .io_in_psum(PE_Array_8_6_io_in_psum),
    .io_in_flow(PE_Array_8_6_io_in_flow),
    .io_in_shift(PE_Array_8_6_io_in_shift),
    .io_out_activate(PE_Array_8_6_io_out_activate),
    .io_out_weight(PE_Array_8_6_io_out_weight),
    .io_out_psum(PE_Array_8_6_io_out_psum)
  );
  basic_PE PE_Array_8_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_7_clock),
    .reset(PE_Array_8_7_reset),
    .io_in_activate(PE_Array_8_7_io_in_activate),
    .io_in_weight(PE_Array_8_7_io_in_weight),
    .io_in_psum(PE_Array_8_7_io_in_psum),
    .io_in_flow(PE_Array_8_7_io_in_flow),
    .io_in_shift(PE_Array_8_7_io_in_shift),
    .io_out_activate(PE_Array_8_7_io_out_activate),
    .io_out_weight(PE_Array_8_7_io_out_weight),
    .io_out_psum(PE_Array_8_7_io_out_psum)
  );
  basic_PE PE_Array_8_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_8_clock),
    .reset(PE_Array_8_8_reset),
    .io_in_activate(PE_Array_8_8_io_in_activate),
    .io_in_weight(PE_Array_8_8_io_in_weight),
    .io_in_psum(PE_Array_8_8_io_in_psum),
    .io_in_flow(PE_Array_8_8_io_in_flow),
    .io_in_shift(PE_Array_8_8_io_in_shift),
    .io_out_activate(PE_Array_8_8_io_out_activate),
    .io_out_weight(PE_Array_8_8_io_out_weight),
    .io_out_psum(PE_Array_8_8_io_out_psum)
  );
  basic_PE PE_Array_8_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_9_clock),
    .reset(PE_Array_8_9_reset),
    .io_in_activate(PE_Array_8_9_io_in_activate),
    .io_in_weight(PE_Array_8_9_io_in_weight),
    .io_in_psum(PE_Array_8_9_io_in_psum),
    .io_in_flow(PE_Array_8_9_io_in_flow),
    .io_in_shift(PE_Array_8_9_io_in_shift),
    .io_out_activate(PE_Array_8_9_io_out_activate),
    .io_out_weight(PE_Array_8_9_io_out_weight),
    .io_out_psum(PE_Array_8_9_io_out_psum)
  );
  basic_PE PE_Array_8_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_10_clock),
    .reset(PE_Array_8_10_reset),
    .io_in_activate(PE_Array_8_10_io_in_activate),
    .io_in_weight(PE_Array_8_10_io_in_weight),
    .io_in_psum(PE_Array_8_10_io_in_psum),
    .io_in_flow(PE_Array_8_10_io_in_flow),
    .io_in_shift(PE_Array_8_10_io_in_shift),
    .io_out_activate(PE_Array_8_10_io_out_activate),
    .io_out_weight(PE_Array_8_10_io_out_weight),
    .io_out_psum(PE_Array_8_10_io_out_psum)
  );
  basic_PE PE_Array_8_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_11_clock),
    .reset(PE_Array_8_11_reset),
    .io_in_activate(PE_Array_8_11_io_in_activate),
    .io_in_weight(PE_Array_8_11_io_in_weight),
    .io_in_psum(PE_Array_8_11_io_in_psum),
    .io_in_flow(PE_Array_8_11_io_in_flow),
    .io_in_shift(PE_Array_8_11_io_in_shift),
    .io_out_activate(PE_Array_8_11_io_out_activate),
    .io_out_weight(PE_Array_8_11_io_out_weight),
    .io_out_psum(PE_Array_8_11_io_out_psum)
  );
  basic_PE PE_Array_8_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_12_clock),
    .reset(PE_Array_8_12_reset),
    .io_in_activate(PE_Array_8_12_io_in_activate),
    .io_in_weight(PE_Array_8_12_io_in_weight),
    .io_in_psum(PE_Array_8_12_io_in_psum),
    .io_in_flow(PE_Array_8_12_io_in_flow),
    .io_in_shift(PE_Array_8_12_io_in_shift),
    .io_out_activate(PE_Array_8_12_io_out_activate),
    .io_out_weight(PE_Array_8_12_io_out_weight),
    .io_out_psum(PE_Array_8_12_io_out_psum)
  );
  basic_PE PE_Array_8_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_13_clock),
    .reset(PE_Array_8_13_reset),
    .io_in_activate(PE_Array_8_13_io_in_activate),
    .io_in_weight(PE_Array_8_13_io_in_weight),
    .io_in_psum(PE_Array_8_13_io_in_psum),
    .io_in_flow(PE_Array_8_13_io_in_flow),
    .io_in_shift(PE_Array_8_13_io_in_shift),
    .io_out_activate(PE_Array_8_13_io_out_activate),
    .io_out_weight(PE_Array_8_13_io_out_weight),
    .io_out_psum(PE_Array_8_13_io_out_psum)
  );
  basic_PE PE_Array_8_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_14_clock),
    .reset(PE_Array_8_14_reset),
    .io_in_activate(PE_Array_8_14_io_in_activate),
    .io_in_weight(PE_Array_8_14_io_in_weight),
    .io_in_psum(PE_Array_8_14_io_in_psum),
    .io_in_flow(PE_Array_8_14_io_in_flow),
    .io_in_shift(PE_Array_8_14_io_in_shift),
    .io_out_activate(PE_Array_8_14_io_out_activate),
    .io_out_weight(PE_Array_8_14_io_out_weight),
    .io_out_psum(PE_Array_8_14_io_out_psum)
  );
  basic_PE PE_Array_8_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_15_clock),
    .reset(PE_Array_8_15_reset),
    .io_in_activate(PE_Array_8_15_io_in_activate),
    .io_in_weight(PE_Array_8_15_io_in_weight),
    .io_in_psum(PE_Array_8_15_io_in_psum),
    .io_in_flow(PE_Array_8_15_io_in_flow),
    .io_in_shift(PE_Array_8_15_io_in_shift),
    .io_out_activate(PE_Array_8_15_io_out_activate),
    .io_out_weight(PE_Array_8_15_io_out_weight),
    .io_out_psum(PE_Array_8_15_io_out_psum)
  );
  basic_PE PE_Array_9_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_0_clock),
    .reset(PE_Array_9_0_reset),
    .io_in_activate(PE_Array_9_0_io_in_activate),
    .io_in_weight(PE_Array_9_0_io_in_weight),
    .io_in_psum(PE_Array_9_0_io_in_psum),
    .io_in_flow(PE_Array_9_0_io_in_flow),
    .io_in_shift(PE_Array_9_0_io_in_shift),
    .io_out_activate(PE_Array_9_0_io_out_activate),
    .io_out_weight(PE_Array_9_0_io_out_weight),
    .io_out_psum(PE_Array_9_0_io_out_psum)
  );
  basic_PE PE_Array_9_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_1_clock),
    .reset(PE_Array_9_1_reset),
    .io_in_activate(PE_Array_9_1_io_in_activate),
    .io_in_weight(PE_Array_9_1_io_in_weight),
    .io_in_psum(PE_Array_9_1_io_in_psum),
    .io_in_flow(PE_Array_9_1_io_in_flow),
    .io_in_shift(PE_Array_9_1_io_in_shift),
    .io_out_activate(PE_Array_9_1_io_out_activate),
    .io_out_weight(PE_Array_9_1_io_out_weight),
    .io_out_psum(PE_Array_9_1_io_out_psum)
  );
  basic_PE PE_Array_9_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_2_clock),
    .reset(PE_Array_9_2_reset),
    .io_in_activate(PE_Array_9_2_io_in_activate),
    .io_in_weight(PE_Array_9_2_io_in_weight),
    .io_in_psum(PE_Array_9_2_io_in_psum),
    .io_in_flow(PE_Array_9_2_io_in_flow),
    .io_in_shift(PE_Array_9_2_io_in_shift),
    .io_out_activate(PE_Array_9_2_io_out_activate),
    .io_out_weight(PE_Array_9_2_io_out_weight),
    .io_out_psum(PE_Array_9_2_io_out_psum)
  );
  basic_PE PE_Array_9_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_3_clock),
    .reset(PE_Array_9_3_reset),
    .io_in_activate(PE_Array_9_3_io_in_activate),
    .io_in_weight(PE_Array_9_3_io_in_weight),
    .io_in_psum(PE_Array_9_3_io_in_psum),
    .io_in_flow(PE_Array_9_3_io_in_flow),
    .io_in_shift(PE_Array_9_3_io_in_shift),
    .io_out_activate(PE_Array_9_3_io_out_activate),
    .io_out_weight(PE_Array_9_3_io_out_weight),
    .io_out_psum(PE_Array_9_3_io_out_psum)
  );
  basic_PE PE_Array_9_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_4_clock),
    .reset(PE_Array_9_4_reset),
    .io_in_activate(PE_Array_9_4_io_in_activate),
    .io_in_weight(PE_Array_9_4_io_in_weight),
    .io_in_psum(PE_Array_9_4_io_in_psum),
    .io_in_flow(PE_Array_9_4_io_in_flow),
    .io_in_shift(PE_Array_9_4_io_in_shift),
    .io_out_activate(PE_Array_9_4_io_out_activate),
    .io_out_weight(PE_Array_9_4_io_out_weight),
    .io_out_psum(PE_Array_9_4_io_out_psum)
  );
  basic_PE PE_Array_9_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_5_clock),
    .reset(PE_Array_9_5_reset),
    .io_in_activate(PE_Array_9_5_io_in_activate),
    .io_in_weight(PE_Array_9_5_io_in_weight),
    .io_in_psum(PE_Array_9_5_io_in_psum),
    .io_in_flow(PE_Array_9_5_io_in_flow),
    .io_in_shift(PE_Array_9_5_io_in_shift),
    .io_out_activate(PE_Array_9_5_io_out_activate),
    .io_out_weight(PE_Array_9_5_io_out_weight),
    .io_out_psum(PE_Array_9_5_io_out_psum)
  );
  basic_PE PE_Array_9_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_6_clock),
    .reset(PE_Array_9_6_reset),
    .io_in_activate(PE_Array_9_6_io_in_activate),
    .io_in_weight(PE_Array_9_6_io_in_weight),
    .io_in_psum(PE_Array_9_6_io_in_psum),
    .io_in_flow(PE_Array_9_6_io_in_flow),
    .io_in_shift(PE_Array_9_6_io_in_shift),
    .io_out_activate(PE_Array_9_6_io_out_activate),
    .io_out_weight(PE_Array_9_6_io_out_weight),
    .io_out_psum(PE_Array_9_6_io_out_psum)
  );
  basic_PE PE_Array_9_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_7_clock),
    .reset(PE_Array_9_7_reset),
    .io_in_activate(PE_Array_9_7_io_in_activate),
    .io_in_weight(PE_Array_9_7_io_in_weight),
    .io_in_psum(PE_Array_9_7_io_in_psum),
    .io_in_flow(PE_Array_9_7_io_in_flow),
    .io_in_shift(PE_Array_9_7_io_in_shift),
    .io_out_activate(PE_Array_9_7_io_out_activate),
    .io_out_weight(PE_Array_9_7_io_out_weight),
    .io_out_psum(PE_Array_9_7_io_out_psum)
  );
  basic_PE PE_Array_9_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_8_clock),
    .reset(PE_Array_9_8_reset),
    .io_in_activate(PE_Array_9_8_io_in_activate),
    .io_in_weight(PE_Array_9_8_io_in_weight),
    .io_in_psum(PE_Array_9_8_io_in_psum),
    .io_in_flow(PE_Array_9_8_io_in_flow),
    .io_in_shift(PE_Array_9_8_io_in_shift),
    .io_out_activate(PE_Array_9_8_io_out_activate),
    .io_out_weight(PE_Array_9_8_io_out_weight),
    .io_out_psum(PE_Array_9_8_io_out_psum)
  );
  basic_PE PE_Array_9_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_9_clock),
    .reset(PE_Array_9_9_reset),
    .io_in_activate(PE_Array_9_9_io_in_activate),
    .io_in_weight(PE_Array_9_9_io_in_weight),
    .io_in_psum(PE_Array_9_9_io_in_psum),
    .io_in_flow(PE_Array_9_9_io_in_flow),
    .io_in_shift(PE_Array_9_9_io_in_shift),
    .io_out_activate(PE_Array_9_9_io_out_activate),
    .io_out_weight(PE_Array_9_9_io_out_weight),
    .io_out_psum(PE_Array_9_9_io_out_psum)
  );
  basic_PE PE_Array_9_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_10_clock),
    .reset(PE_Array_9_10_reset),
    .io_in_activate(PE_Array_9_10_io_in_activate),
    .io_in_weight(PE_Array_9_10_io_in_weight),
    .io_in_psum(PE_Array_9_10_io_in_psum),
    .io_in_flow(PE_Array_9_10_io_in_flow),
    .io_in_shift(PE_Array_9_10_io_in_shift),
    .io_out_activate(PE_Array_9_10_io_out_activate),
    .io_out_weight(PE_Array_9_10_io_out_weight),
    .io_out_psum(PE_Array_9_10_io_out_psum)
  );
  basic_PE PE_Array_9_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_11_clock),
    .reset(PE_Array_9_11_reset),
    .io_in_activate(PE_Array_9_11_io_in_activate),
    .io_in_weight(PE_Array_9_11_io_in_weight),
    .io_in_psum(PE_Array_9_11_io_in_psum),
    .io_in_flow(PE_Array_9_11_io_in_flow),
    .io_in_shift(PE_Array_9_11_io_in_shift),
    .io_out_activate(PE_Array_9_11_io_out_activate),
    .io_out_weight(PE_Array_9_11_io_out_weight),
    .io_out_psum(PE_Array_9_11_io_out_psum)
  );
  basic_PE PE_Array_9_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_12_clock),
    .reset(PE_Array_9_12_reset),
    .io_in_activate(PE_Array_9_12_io_in_activate),
    .io_in_weight(PE_Array_9_12_io_in_weight),
    .io_in_psum(PE_Array_9_12_io_in_psum),
    .io_in_flow(PE_Array_9_12_io_in_flow),
    .io_in_shift(PE_Array_9_12_io_in_shift),
    .io_out_activate(PE_Array_9_12_io_out_activate),
    .io_out_weight(PE_Array_9_12_io_out_weight),
    .io_out_psum(PE_Array_9_12_io_out_psum)
  );
  basic_PE PE_Array_9_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_13_clock),
    .reset(PE_Array_9_13_reset),
    .io_in_activate(PE_Array_9_13_io_in_activate),
    .io_in_weight(PE_Array_9_13_io_in_weight),
    .io_in_psum(PE_Array_9_13_io_in_psum),
    .io_in_flow(PE_Array_9_13_io_in_flow),
    .io_in_shift(PE_Array_9_13_io_in_shift),
    .io_out_activate(PE_Array_9_13_io_out_activate),
    .io_out_weight(PE_Array_9_13_io_out_weight),
    .io_out_psum(PE_Array_9_13_io_out_psum)
  );
  basic_PE PE_Array_9_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_14_clock),
    .reset(PE_Array_9_14_reset),
    .io_in_activate(PE_Array_9_14_io_in_activate),
    .io_in_weight(PE_Array_9_14_io_in_weight),
    .io_in_psum(PE_Array_9_14_io_in_psum),
    .io_in_flow(PE_Array_9_14_io_in_flow),
    .io_in_shift(PE_Array_9_14_io_in_shift),
    .io_out_activate(PE_Array_9_14_io_out_activate),
    .io_out_weight(PE_Array_9_14_io_out_weight),
    .io_out_psum(PE_Array_9_14_io_out_psum)
  );
  basic_PE PE_Array_9_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_15_clock),
    .reset(PE_Array_9_15_reset),
    .io_in_activate(PE_Array_9_15_io_in_activate),
    .io_in_weight(PE_Array_9_15_io_in_weight),
    .io_in_psum(PE_Array_9_15_io_in_psum),
    .io_in_flow(PE_Array_9_15_io_in_flow),
    .io_in_shift(PE_Array_9_15_io_in_shift),
    .io_out_activate(PE_Array_9_15_io_out_activate),
    .io_out_weight(PE_Array_9_15_io_out_weight),
    .io_out_psum(PE_Array_9_15_io_out_psum)
  );
  basic_PE PE_Array_10_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_0_clock),
    .reset(PE_Array_10_0_reset),
    .io_in_activate(PE_Array_10_0_io_in_activate),
    .io_in_weight(PE_Array_10_0_io_in_weight),
    .io_in_psum(PE_Array_10_0_io_in_psum),
    .io_in_flow(PE_Array_10_0_io_in_flow),
    .io_in_shift(PE_Array_10_0_io_in_shift),
    .io_out_activate(PE_Array_10_0_io_out_activate),
    .io_out_weight(PE_Array_10_0_io_out_weight),
    .io_out_psum(PE_Array_10_0_io_out_psum)
  );
  basic_PE PE_Array_10_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_1_clock),
    .reset(PE_Array_10_1_reset),
    .io_in_activate(PE_Array_10_1_io_in_activate),
    .io_in_weight(PE_Array_10_1_io_in_weight),
    .io_in_psum(PE_Array_10_1_io_in_psum),
    .io_in_flow(PE_Array_10_1_io_in_flow),
    .io_in_shift(PE_Array_10_1_io_in_shift),
    .io_out_activate(PE_Array_10_1_io_out_activate),
    .io_out_weight(PE_Array_10_1_io_out_weight),
    .io_out_psum(PE_Array_10_1_io_out_psum)
  );
  basic_PE PE_Array_10_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_2_clock),
    .reset(PE_Array_10_2_reset),
    .io_in_activate(PE_Array_10_2_io_in_activate),
    .io_in_weight(PE_Array_10_2_io_in_weight),
    .io_in_psum(PE_Array_10_2_io_in_psum),
    .io_in_flow(PE_Array_10_2_io_in_flow),
    .io_in_shift(PE_Array_10_2_io_in_shift),
    .io_out_activate(PE_Array_10_2_io_out_activate),
    .io_out_weight(PE_Array_10_2_io_out_weight),
    .io_out_psum(PE_Array_10_2_io_out_psum)
  );
  basic_PE PE_Array_10_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_3_clock),
    .reset(PE_Array_10_3_reset),
    .io_in_activate(PE_Array_10_3_io_in_activate),
    .io_in_weight(PE_Array_10_3_io_in_weight),
    .io_in_psum(PE_Array_10_3_io_in_psum),
    .io_in_flow(PE_Array_10_3_io_in_flow),
    .io_in_shift(PE_Array_10_3_io_in_shift),
    .io_out_activate(PE_Array_10_3_io_out_activate),
    .io_out_weight(PE_Array_10_3_io_out_weight),
    .io_out_psum(PE_Array_10_3_io_out_psum)
  );
  basic_PE PE_Array_10_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_4_clock),
    .reset(PE_Array_10_4_reset),
    .io_in_activate(PE_Array_10_4_io_in_activate),
    .io_in_weight(PE_Array_10_4_io_in_weight),
    .io_in_psum(PE_Array_10_4_io_in_psum),
    .io_in_flow(PE_Array_10_4_io_in_flow),
    .io_in_shift(PE_Array_10_4_io_in_shift),
    .io_out_activate(PE_Array_10_4_io_out_activate),
    .io_out_weight(PE_Array_10_4_io_out_weight),
    .io_out_psum(PE_Array_10_4_io_out_psum)
  );
  basic_PE PE_Array_10_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_5_clock),
    .reset(PE_Array_10_5_reset),
    .io_in_activate(PE_Array_10_5_io_in_activate),
    .io_in_weight(PE_Array_10_5_io_in_weight),
    .io_in_psum(PE_Array_10_5_io_in_psum),
    .io_in_flow(PE_Array_10_5_io_in_flow),
    .io_in_shift(PE_Array_10_5_io_in_shift),
    .io_out_activate(PE_Array_10_5_io_out_activate),
    .io_out_weight(PE_Array_10_5_io_out_weight),
    .io_out_psum(PE_Array_10_5_io_out_psum)
  );
  basic_PE PE_Array_10_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_6_clock),
    .reset(PE_Array_10_6_reset),
    .io_in_activate(PE_Array_10_6_io_in_activate),
    .io_in_weight(PE_Array_10_6_io_in_weight),
    .io_in_psum(PE_Array_10_6_io_in_psum),
    .io_in_flow(PE_Array_10_6_io_in_flow),
    .io_in_shift(PE_Array_10_6_io_in_shift),
    .io_out_activate(PE_Array_10_6_io_out_activate),
    .io_out_weight(PE_Array_10_6_io_out_weight),
    .io_out_psum(PE_Array_10_6_io_out_psum)
  );
  basic_PE PE_Array_10_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_7_clock),
    .reset(PE_Array_10_7_reset),
    .io_in_activate(PE_Array_10_7_io_in_activate),
    .io_in_weight(PE_Array_10_7_io_in_weight),
    .io_in_psum(PE_Array_10_7_io_in_psum),
    .io_in_flow(PE_Array_10_7_io_in_flow),
    .io_in_shift(PE_Array_10_7_io_in_shift),
    .io_out_activate(PE_Array_10_7_io_out_activate),
    .io_out_weight(PE_Array_10_7_io_out_weight),
    .io_out_psum(PE_Array_10_7_io_out_psum)
  );
  basic_PE PE_Array_10_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_8_clock),
    .reset(PE_Array_10_8_reset),
    .io_in_activate(PE_Array_10_8_io_in_activate),
    .io_in_weight(PE_Array_10_8_io_in_weight),
    .io_in_psum(PE_Array_10_8_io_in_psum),
    .io_in_flow(PE_Array_10_8_io_in_flow),
    .io_in_shift(PE_Array_10_8_io_in_shift),
    .io_out_activate(PE_Array_10_8_io_out_activate),
    .io_out_weight(PE_Array_10_8_io_out_weight),
    .io_out_psum(PE_Array_10_8_io_out_psum)
  );
  basic_PE PE_Array_10_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_9_clock),
    .reset(PE_Array_10_9_reset),
    .io_in_activate(PE_Array_10_9_io_in_activate),
    .io_in_weight(PE_Array_10_9_io_in_weight),
    .io_in_psum(PE_Array_10_9_io_in_psum),
    .io_in_flow(PE_Array_10_9_io_in_flow),
    .io_in_shift(PE_Array_10_9_io_in_shift),
    .io_out_activate(PE_Array_10_9_io_out_activate),
    .io_out_weight(PE_Array_10_9_io_out_weight),
    .io_out_psum(PE_Array_10_9_io_out_psum)
  );
  basic_PE PE_Array_10_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_10_clock),
    .reset(PE_Array_10_10_reset),
    .io_in_activate(PE_Array_10_10_io_in_activate),
    .io_in_weight(PE_Array_10_10_io_in_weight),
    .io_in_psum(PE_Array_10_10_io_in_psum),
    .io_in_flow(PE_Array_10_10_io_in_flow),
    .io_in_shift(PE_Array_10_10_io_in_shift),
    .io_out_activate(PE_Array_10_10_io_out_activate),
    .io_out_weight(PE_Array_10_10_io_out_weight),
    .io_out_psum(PE_Array_10_10_io_out_psum)
  );
  basic_PE PE_Array_10_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_11_clock),
    .reset(PE_Array_10_11_reset),
    .io_in_activate(PE_Array_10_11_io_in_activate),
    .io_in_weight(PE_Array_10_11_io_in_weight),
    .io_in_psum(PE_Array_10_11_io_in_psum),
    .io_in_flow(PE_Array_10_11_io_in_flow),
    .io_in_shift(PE_Array_10_11_io_in_shift),
    .io_out_activate(PE_Array_10_11_io_out_activate),
    .io_out_weight(PE_Array_10_11_io_out_weight),
    .io_out_psum(PE_Array_10_11_io_out_psum)
  );
  basic_PE PE_Array_10_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_12_clock),
    .reset(PE_Array_10_12_reset),
    .io_in_activate(PE_Array_10_12_io_in_activate),
    .io_in_weight(PE_Array_10_12_io_in_weight),
    .io_in_psum(PE_Array_10_12_io_in_psum),
    .io_in_flow(PE_Array_10_12_io_in_flow),
    .io_in_shift(PE_Array_10_12_io_in_shift),
    .io_out_activate(PE_Array_10_12_io_out_activate),
    .io_out_weight(PE_Array_10_12_io_out_weight),
    .io_out_psum(PE_Array_10_12_io_out_psum)
  );
  basic_PE PE_Array_10_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_13_clock),
    .reset(PE_Array_10_13_reset),
    .io_in_activate(PE_Array_10_13_io_in_activate),
    .io_in_weight(PE_Array_10_13_io_in_weight),
    .io_in_psum(PE_Array_10_13_io_in_psum),
    .io_in_flow(PE_Array_10_13_io_in_flow),
    .io_in_shift(PE_Array_10_13_io_in_shift),
    .io_out_activate(PE_Array_10_13_io_out_activate),
    .io_out_weight(PE_Array_10_13_io_out_weight),
    .io_out_psum(PE_Array_10_13_io_out_psum)
  );
  basic_PE PE_Array_10_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_14_clock),
    .reset(PE_Array_10_14_reset),
    .io_in_activate(PE_Array_10_14_io_in_activate),
    .io_in_weight(PE_Array_10_14_io_in_weight),
    .io_in_psum(PE_Array_10_14_io_in_psum),
    .io_in_flow(PE_Array_10_14_io_in_flow),
    .io_in_shift(PE_Array_10_14_io_in_shift),
    .io_out_activate(PE_Array_10_14_io_out_activate),
    .io_out_weight(PE_Array_10_14_io_out_weight),
    .io_out_psum(PE_Array_10_14_io_out_psum)
  );
  basic_PE PE_Array_10_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_15_clock),
    .reset(PE_Array_10_15_reset),
    .io_in_activate(PE_Array_10_15_io_in_activate),
    .io_in_weight(PE_Array_10_15_io_in_weight),
    .io_in_psum(PE_Array_10_15_io_in_psum),
    .io_in_flow(PE_Array_10_15_io_in_flow),
    .io_in_shift(PE_Array_10_15_io_in_shift),
    .io_out_activate(PE_Array_10_15_io_out_activate),
    .io_out_weight(PE_Array_10_15_io_out_weight),
    .io_out_psum(PE_Array_10_15_io_out_psum)
  );
  basic_PE PE_Array_11_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_0_clock),
    .reset(PE_Array_11_0_reset),
    .io_in_activate(PE_Array_11_0_io_in_activate),
    .io_in_weight(PE_Array_11_0_io_in_weight),
    .io_in_psum(PE_Array_11_0_io_in_psum),
    .io_in_flow(PE_Array_11_0_io_in_flow),
    .io_in_shift(PE_Array_11_0_io_in_shift),
    .io_out_activate(PE_Array_11_0_io_out_activate),
    .io_out_weight(PE_Array_11_0_io_out_weight),
    .io_out_psum(PE_Array_11_0_io_out_psum)
  );
  basic_PE PE_Array_11_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_1_clock),
    .reset(PE_Array_11_1_reset),
    .io_in_activate(PE_Array_11_1_io_in_activate),
    .io_in_weight(PE_Array_11_1_io_in_weight),
    .io_in_psum(PE_Array_11_1_io_in_psum),
    .io_in_flow(PE_Array_11_1_io_in_flow),
    .io_in_shift(PE_Array_11_1_io_in_shift),
    .io_out_activate(PE_Array_11_1_io_out_activate),
    .io_out_weight(PE_Array_11_1_io_out_weight),
    .io_out_psum(PE_Array_11_1_io_out_psum)
  );
  basic_PE PE_Array_11_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_2_clock),
    .reset(PE_Array_11_2_reset),
    .io_in_activate(PE_Array_11_2_io_in_activate),
    .io_in_weight(PE_Array_11_2_io_in_weight),
    .io_in_psum(PE_Array_11_2_io_in_psum),
    .io_in_flow(PE_Array_11_2_io_in_flow),
    .io_in_shift(PE_Array_11_2_io_in_shift),
    .io_out_activate(PE_Array_11_2_io_out_activate),
    .io_out_weight(PE_Array_11_2_io_out_weight),
    .io_out_psum(PE_Array_11_2_io_out_psum)
  );
  basic_PE PE_Array_11_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_3_clock),
    .reset(PE_Array_11_3_reset),
    .io_in_activate(PE_Array_11_3_io_in_activate),
    .io_in_weight(PE_Array_11_3_io_in_weight),
    .io_in_psum(PE_Array_11_3_io_in_psum),
    .io_in_flow(PE_Array_11_3_io_in_flow),
    .io_in_shift(PE_Array_11_3_io_in_shift),
    .io_out_activate(PE_Array_11_3_io_out_activate),
    .io_out_weight(PE_Array_11_3_io_out_weight),
    .io_out_psum(PE_Array_11_3_io_out_psum)
  );
  basic_PE PE_Array_11_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_4_clock),
    .reset(PE_Array_11_4_reset),
    .io_in_activate(PE_Array_11_4_io_in_activate),
    .io_in_weight(PE_Array_11_4_io_in_weight),
    .io_in_psum(PE_Array_11_4_io_in_psum),
    .io_in_flow(PE_Array_11_4_io_in_flow),
    .io_in_shift(PE_Array_11_4_io_in_shift),
    .io_out_activate(PE_Array_11_4_io_out_activate),
    .io_out_weight(PE_Array_11_4_io_out_weight),
    .io_out_psum(PE_Array_11_4_io_out_psum)
  );
  basic_PE PE_Array_11_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_5_clock),
    .reset(PE_Array_11_5_reset),
    .io_in_activate(PE_Array_11_5_io_in_activate),
    .io_in_weight(PE_Array_11_5_io_in_weight),
    .io_in_psum(PE_Array_11_5_io_in_psum),
    .io_in_flow(PE_Array_11_5_io_in_flow),
    .io_in_shift(PE_Array_11_5_io_in_shift),
    .io_out_activate(PE_Array_11_5_io_out_activate),
    .io_out_weight(PE_Array_11_5_io_out_weight),
    .io_out_psum(PE_Array_11_5_io_out_psum)
  );
  basic_PE PE_Array_11_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_6_clock),
    .reset(PE_Array_11_6_reset),
    .io_in_activate(PE_Array_11_6_io_in_activate),
    .io_in_weight(PE_Array_11_6_io_in_weight),
    .io_in_psum(PE_Array_11_6_io_in_psum),
    .io_in_flow(PE_Array_11_6_io_in_flow),
    .io_in_shift(PE_Array_11_6_io_in_shift),
    .io_out_activate(PE_Array_11_6_io_out_activate),
    .io_out_weight(PE_Array_11_6_io_out_weight),
    .io_out_psum(PE_Array_11_6_io_out_psum)
  );
  basic_PE PE_Array_11_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_7_clock),
    .reset(PE_Array_11_7_reset),
    .io_in_activate(PE_Array_11_7_io_in_activate),
    .io_in_weight(PE_Array_11_7_io_in_weight),
    .io_in_psum(PE_Array_11_7_io_in_psum),
    .io_in_flow(PE_Array_11_7_io_in_flow),
    .io_in_shift(PE_Array_11_7_io_in_shift),
    .io_out_activate(PE_Array_11_7_io_out_activate),
    .io_out_weight(PE_Array_11_7_io_out_weight),
    .io_out_psum(PE_Array_11_7_io_out_psum)
  );
  basic_PE PE_Array_11_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_8_clock),
    .reset(PE_Array_11_8_reset),
    .io_in_activate(PE_Array_11_8_io_in_activate),
    .io_in_weight(PE_Array_11_8_io_in_weight),
    .io_in_psum(PE_Array_11_8_io_in_psum),
    .io_in_flow(PE_Array_11_8_io_in_flow),
    .io_in_shift(PE_Array_11_8_io_in_shift),
    .io_out_activate(PE_Array_11_8_io_out_activate),
    .io_out_weight(PE_Array_11_8_io_out_weight),
    .io_out_psum(PE_Array_11_8_io_out_psum)
  );
  basic_PE PE_Array_11_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_9_clock),
    .reset(PE_Array_11_9_reset),
    .io_in_activate(PE_Array_11_9_io_in_activate),
    .io_in_weight(PE_Array_11_9_io_in_weight),
    .io_in_psum(PE_Array_11_9_io_in_psum),
    .io_in_flow(PE_Array_11_9_io_in_flow),
    .io_in_shift(PE_Array_11_9_io_in_shift),
    .io_out_activate(PE_Array_11_9_io_out_activate),
    .io_out_weight(PE_Array_11_9_io_out_weight),
    .io_out_psum(PE_Array_11_9_io_out_psum)
  );
  basic_PE PE_Array_11_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_10_clock),
    .reset(PE_Array_11_10_reset),
    .io_in_activate(PE_Array_11_10_io_in_activate),
    .io_in_weight(PE_Array_11_10_io_in_weight),
    .io_in_psum(PE_Array_11_10_io_in_psum),
    .io_in_flow(PE_Array_11_10_io_in_flow),
    .io_in_shift(PE_Array_11_10_io_in_shift),
    .io_out_activate(PE_Array_11_10_io_out_activate),
    .io_out_weight(PE_Array_11_10_io_out_weight),
    .io_out_psum(PE_Array_11_10_io_out_psum)
  );
  basic_PE PE_Array_11_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_11_clock),
    .reset(PE_Array_11_11_reset),
    .io_in_activate(PE_Array_11_11_io_in_activate),
    .io_in_weight(PE_Array_11_11_io_in_weight),
    .io_in_psum(PE_Array_11_11_io_in_psum),
    .io_in_flow(PE_Array_11_11_io_in_flow),
    .io_in_shift(PE_Array_11_11_io_in_shift),
    .io_out_activate(PE_Array_11_11_io_out_activate),
    .io_out_weight(PE_Array_11_11_io_out_weight),
    .io_out_psum(PE_Array_11_11_io_out_psum)
  );
  basic_PE PE_Array_11_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_12_clock),
    .reset(PE_Array_11_12_reset),
    .io_in_activate(PE_Array_11_12_io_in_activate),
    .io_in_weight(PE_Array_11_12_io_in_weight),
    .io_in_psum(PE_Array_11_12_io_in_psum),
    .io_in_flow(PE_Array_11_12_io_in_flow),
    .io_in_shift(PE_Array_11_12_io_in_shift),
    .io_out_activate(PE_Array_11_12_io_out_activate),
    .io_out_weight(PE_Array_11_12_io_out_weight),
    .io_out_psum(PE_Array_11_12_io_out_psum)
  );
  basic_PE PE_Array_11_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_13_clock),
    .reset(PE_Array_11_13_reset),
    .io_in_activate(PE_Array_11_13_io_in_activate),
    .io_in_weight(PE_Array_11_13_io_in_weight),
    .io_in_psum(PE_Array_11_13_io_in_psum),
    .io_in_flow(PE_Array_11_13_io_in_flow),
    .io_in_shift(PE_Array_11_13_io_in_shift),
    .io_out_activate(PE_Array_11_13_io_out_activate),
    .io_out_weight(PE_Array_11_13_io_out_weight),
    .io_out_psum(PE_Array_11_13_io_out_psum)
  );
  basic_PE PE_Array_11_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_14_clock),
    .reset(PE_Array_11_14_reset),
    .io_in_activate(PE_Array_11_14_io_in_activate),
    .io_in_weight(PE_Array_11_14_io_in_weight),
    .io_in_psum(PE_Array_11_14_io_in_psum),
    .io_in_flow(PE_Array_11_14_io_in_flow),
    .io_in_shift(PE_Array_11_14_io_in_shift),
    .io_out_activate(PE_Array_11_14_io_out_activate),
    .io_out_weight(PE_Array_11_14_io_out_weight),
    .io_out_psum(PE_Array_11_14_io_out_psum)
  );
  basic_PE PE_Array_11_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_15_clock),
    .reset(PE_Array_11_15_reset),
    .io_in_activate(PE_Array_11_15_io_in_activate),
    .io_in_weight(PE_Array_11_15_io_in_weight),
    .io_in_psum(PE_Array_11_15_io_in_psum),
    .io_in_flow(PE_Array_11_15_io_in_flow),
    .io_in_shift(PE_Array_11_15_io_in_shift),
    .io_out_activate(PE_Array_11_15_io_out_activate),
    .io_out_weight(PE_Array_11_15_io_out_weight),
    .io_out_psum(PE_Array_11_15_io_out_psum)
  );
  basic_PE PE_Array_12_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_0_clock),
    .reset(PE_Array_12_0_reset),
    .io_in_activate(PE_Array_12_0_io_in_activate),
    .io_in_weight(PE_Array_12_0_io_in_weight),
    .io_in_psum(PE_Array_12_0_io_in_psum),
    .io_in_flow(PE_Array_12_0_io_in_flow),
    .io_in_shift(PE_Array_12_0_io_in_shift),
    .io_out_activate(PE_Array_12_0_io_out_activate),
    .io_out_weight(PE_Array_12_0_io_out_weight),
    .io_out_psum(PE_Array_12_0_io_out_psum)
  );
  basic_PE PE_Array_12_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_1_clock),
    .reset(PE_Array_12_1_reset),
    .io_in_activate(PE_Array_12_1_io_in_activate),
    .io_in_weight(PE_Array_12_1_io_in_weight),
    .io_in_psum(PE_Array_12_1_io_in_psum),
    .io_in_flow(PE_Array_12_1_io_in_flow),
    .io_in_shift(PE_Array_12_1_io_in_shift),
    .io_out_activate(PE_Array_12_1_io_out_activate),
    .io_out_weight(PE_Array_12_1_io_out_weight),
    .io_out_psum(PE_Array_12_1_io_out_psum)
  );
  basic_PE PE_Array_12_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_2_clock),
    .reset(PE_Array_12_2_reset),
    .io_in_activate(PE_Array_12_2_io_in_activate),
    .io_in_weight(PE_Array_12_2_io_in_weight),
    .io_in_psum(PE_Array_12_2_io_in_psum),
    .io_in_flow(PE_Array_12_2_io_in_flow),
    .io_in_shift(PE_Array_12_2_io_in_shift),
    .io_out_activate(PE_Array_12_2_io_out_activate),
    .io_out_weight(PE_Array_12_2_io_out_weight),
    .io_out_psum(PE_Array_12_2_io_out_psum)
  );
  basic_PE PE_Array_12_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_3_clock),
    .reset(PE_Array_12_3_reset),
    .io_in_activate(PE_Array_12_3_io_in_activate),
    .io_in_weight(PE_Array_12_3_io_in_weight),
    .io_in_psum(PE_Array_12_3_io_in_psum),
    .io_in_flow(PE_Array_12_3_io_in_flow),
    .io_in_shift(PE_Array_12_3_io_in_shift),
    .io_out_activate(PE_Array_12_3_io_out_activate),
    .io_out_weight(PE_Array_12_3_io_out_weight),
    .io_out_psum(PE_Array_12_3_io_out_psum)
  );
  basic_PE PE_Array_12_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_4_clock),
    .reset(PE_Array_12_4_reset),
    .io_in_activate(PE_Array_12_4_io_in_activate),
    .io_in_weight(PE_Array_12_4_io_in_weight),
    .io_in_psum(PE_Array_12_4_io_in_psum),
    .io_in_flow(PE_Array_12_4_io_in_flow),
    .io_in_shift(PE_Array_12_4_io_in_shift),
    .io_out_activate(PE_Array_12_4_io_out_activate),
    .io_out_weight(PE_Array_12_4_io_out_weight),
    .io_out_psum(PE_Array_12_4_io_out_psum)
  );
  basic_PE PE_Array_12_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_5_clock),
    .reset(PE_Array_12_5_reset),
    .io_in_activate(PE_Array_12_5_io_in_activate),
    .io_in_weight(PE_Array_12_5_io_in_weight),
    .io_in_psum(PE_Array_12_5_io_in_psum),
    .io_in_flow(PE_Array_12_5_io_in_flow),
    .io_in_shift(PE_Array_12_5_io_in_shift),
    .io_out_activate(PE_Array_12_5_io_out_activate),
    .io_out_weight(PE_Array_12_5_io_out_weight),
    .io_out_psum(PE_Array_12_5_io_out_psum)
  );
  basic_PE PE_Array_12_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_6_clock),
    .reset(PE_Array_12_6_reset),
    .io_in_activate(PE_Array_12_6_io_in_activate),
    .io_in_weight(PE_Array_12_6_io_in_weight),
    .io_in_psum(PE_Array_12_6_io_in_psum),
    .io_in_flow(PE_Array_12_6_io_in_flow),
    .io_in_shift(PE_Array_12_6_io_in_shift),
    .io_out_activate(PE_Array_12_6_io_out_activate),
    .io_out_weight(PE_Array_12_6_io_out_weight),
    .io_out_psum(PE_Array_12_6_io_out_psum)
  );
  basic_PE PE_Array_12_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_7_clock),
    .reset(PE_Array_12_7_reset),
    .io_in_activate(PE_Array_12_7_io_in_activate),
    .io_in_weight(PE_Array_12_7_io_in_weight),
    .io_in_psum(PE_Array_12_7_io_in_psum),
    .io_in_flow(PE_Array_12_7_io_in_flow),
    .io_in_shift(PE_Array_12_7_io_in_shift),
    .io_out_activate(PE_Array_12_7_io_out_activate),
    .io_out_weight(PE_Array_12_7_io_out_weight),
    .io_out_psum(PE_Array_12_7_io_out_psum)
  );
  basic_PE PE_Array_12_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_8_clock),
    .reset(PE_Array_12_8_reset),
    .io_in_activate(PE_Array_12_8_io_in_activate),
    .io_in_weight(PE_Array_12_8_io_in_weight),
    .io_in_psum(PE_Array_12_8_io_in_psum),
    .io_in_flow(PE_Array_12_8_io_in_flow),
    .io_in_shift(PE_Array_12_8_io_in_shift),
    .io_out_activate(PE_Array_12_8_io_out_activate),
    .io_out_weight(PE_Array_12_8_io_out_weight),
    .io_out_psum(PE_Array_12_8_io_out_psum)
  );
  basic_PE PE_Array_12_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_9_clock),
    .reset(PE_Array_12_9_reset),
    .io_in_activate(PE_Array_12_9_io_in_activate),
    .io_in_weight(PE_Array_12_9_io_in_weight),
    .io_in_psum(PE_Array_12_9_io_in_psum),
    .io_in_flow(PE_Array_12_9_io_in_flow),
    .io_in_shift(PE_Array_12_9_io_in_shift),
    .io_out_activate(PE_Array_12_9_io_out_activate),
    .io_out_weight(PE_Array_12_9_io_out_weight),
    .io_out_psum(PE_Array_12_9_io_out_psum)
  );
  basic_PE PE_Array_12_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_10_clock),
    .reset(PE_Array_12_10_reset),
    .io_in_activate(PE_Array_12_10_io_in_activate),
    .io_in_weight(PE_Array_12_10_io_in_weight),
    .io_in_psum(PE_Array_12_10_io_in_psum),
    .io_in_flow(PE_Array_12_10_io_in_flow),
    .io_in_shift(PE_Array_12_10_io_in_shift),
    .io_out_activate(PE_Array_12_10_io_out_activate),
    .io_out_weight(PE_Array_12_10_io_out_weight),
    .io_out_psum(PE_Array_12_10_io_out_psum)
  );
  basic_PE PE_Array_12_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_11_clock),
    .reset(PE_Array_12_11_reset),
    .io_in_activate(PE_Array_12_11_io_in_activate),
    .io_in_weight(PE_Array_12_11_io_in_weight),
    .io_in_psum(PE_Array_12_11_io_in_psum),
    .io_in_flow(PE_Array_12_11_io_in_flow),
    .io_in_shift(PE_Array_12_11_io_in_shift),
    .io_out_activate(PE_Array_12_11_io_out_activate),
    .io_out_weight(PE_Array_12_11_io_out_weight),
    .io_out_psum(PE_Array_12_11_io_out_psum)
  );
  basic_PE PE_Array_12_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_12_clock),
    .reset(PE_Array_12_12_reset),
    .io_in_activate(PE_Array_12_12_io_in_activate),
    .io_in_weight(PE_Array_12_12_io_in_weight),
    .io_in_psum(PE_Array_12_12_io_in_psum),
    .io_in_flow(PE_Array_12_12_io_in_flow),
    .io_in_shift(PE_Array_12_12_io_in_shift),
    .io_out_activate(PE_Array_12_12_io_out_activate),
    .io_out_weight(PE_Array_12_12_io_out_weight),
    .io_out_psum(PE_Array_12_12_io_out_psum)
  );
  basic_PE PE_Array_12_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_13_clock),
    .reset(PE_Array_12_13_reset),
    .io_in_activate(PE_Array_12_13_io_in_activate),
    .io_in_weight(PE_Array_12_13_io_in_weight),
    .io_in_psum(PE_Array_12_13_io_in_psum),
    .io_in_flow(PE_Array_12_13_io_in_flow),
    .io_in_shift(PE_Array_12_13_io_in_shift),
    .io_out_activate(PE_Array_12_13_io_out_activate),
    .io_out_weight(PE_Array_12_13_io_out_weight),
    .io_out_psum(PE_Array_12_13_io_out_psum)
  );
  basic_PE PE_Array_12_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_14_clock),
    .reset(PE_Array_12_14_reset),
    .io_in_activate(PE_Array_12_14_io_in_activate),
    .io_in_weight(PE_Array_12_14_io_in_weight),
    .io_in_psum(PE_Array_12_14_io_in_psum),
    .io_in_flow(PE_Array_12_14_io_in_flow),
    .io_in_shift(PE_Array_12_14_io_in_shift),
    .io_out_activate(PE_Array_12_14_io_out_activate),
    .io_out_weight(PE_Array_12_14_io_out_weight),
    .io_out_psum(PE_Array_12_14_io_out_psum)
  );
  basic_PE PE_Array_12_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_15_clock),
    .reset(PE_Array_12_15_reset),
    .io_in_activate(PE_Array_12_15_io_in_activate),
    .io_in_weight(PE_Array_12_15_io_in_weight),
    .io_in_psum(PE_Array_12_15_io_in_psum),
    .io_in_flow(PE_Array_12_15_io_in_flow),
    .io_in_shift(PE_Array_12_15_io_in_shift),
    .io_out_activate(PE_Array_12_15_io_out_activate),
    .io_out_weight(PE_Array_12_15_io_out_weight),
    .io_out_psum(PE_Array_12_15_io_out_psum)
  );
  basic_PE PE_Array_13_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_0_clock),
    .reset(PE_Array_13_0_reset),
    .io_in_activate(PE_Array_13_0_io_in_activate),
    .io_in_weight(PE_Array_13_0_io_in_weight),
    .io_in_psum(PE_Array_13_0_io_in_psum),
    .io_in_flow(PE_Array_13_0_io_in_flow),
    .io_in_shift(PE_Array_13_0_io_in_shift),
    .io_out_activate(PE_Array_13_0_io_out_activate),
    .io_out_weight(PE_Array_13_0_io_out_weight),
    .io_out_psum(PE_Array_13_0_io_out_psum)
  );
  basic_PE PE_Array_13_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_1_clock),
    .reset(PE_Array_13_1_reset),
    .io_in_activate(PE_Array_13_1_io_in_activate),
    .io_in_weight(PE_Array_13_1_io_in_weight),
    .io_in_psum(PE_Array_13_1_io_in_psum),
    .io_in_flow(PE_Array_13_1_io_in_flow),
    .io_in_shift(PE_Array_13_1_io_in_shift),
    .io_out_activate(PE_Array_13_1_io_out_activate),
    .io_out_weight(PE_Array_13_1_io_out_weight),
    .io_out_psum(PE_Array_13_1_io_out_psum)
  );
  basic_PE PE_Array_13_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_2_clock),
    .reset(PE_Array_13_2_reset),
    .io_in_activate(PE_Array_13_2_io_in_activate),
    .io_in_weight(PE_Array_13_2_io_in_weight),
    .io_in_psum(PE_Array_13_2_io_in_psum),
    .io_in_flow(PE_Array_13_2_io_in_flow),
    .io_in_shift(PE_Array_13_2_io_in_shift),
    .io_out_activate(PE_Array_13_2_io_out_activate),
    .io_out_weight(PE_Array_13_2_io_out_weight),
    .io_out_psum(PE_Array_13_2_io_out_psum)
  );
  basic_PE PE_Array_13_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_3_clock),
    .reset(PE_Array_13_3_reset),
    .io_in_activate(PE_Array_13_3_io_in_activate),
    .io_in_weight(PE_Array_13_3_io_in_weight),
    .io_in_psum(PE_Array_13_3_io_in_psum),
    .io_in_flow(PE_Array_13_3_io_in_flow),
    .io_in_shift(PE_Array_13_3_io_in_shift),
    .io_out_activate(PE_Array_13_3_io_out_activate),
    .io_out_weight(PE_Array_13_3_io_out_weight),
    .io_out_psum(PE_Array_13_3_io_out_psum)
  );
  basic_PE PE_Array_13_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_4_clock),
    .reset(PE_Array_13_4_reset),
    .io_in_activate(PE_Array_13_4_io_in_activate),
    .io_in_weight(PE_Array_13_4_io_in_weight),
    .io_in_psum(PE_Array_13_4_io_in_psum),
    .io_in_flow(PE_Array_13_4_io_in_flow),
    .io_in_shift(PE_Array_13_4_io_in_shift),
    .io_out_activate(PE_Array_13_4_io_out_activate),
    .io_out_weight(PE_Array_13_4_io_out_weight),
    .io_out_psum(PE_Array_13_4_io_out_psum)
  );
  basic_PE PE_Array_13_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_5_clock),
    .reset(PE_Array_13_5_reset),
    .io_in_activate(PE_Array_13_5_io_in_activate),
    .io_in_weight(PE_Array_13_5_io_in_weight),
    .io_in_psum(PE_Array_13_5_io_in_psum),
    .io_in_flow(PE_Array_13_5_io_in_flow),
    .io_in_shift(PE_Array_13_5_io_in_shift),
    .io_out_activate(PE_Array_13_5_io_out_activate),
    .io_out_weight(PE_Array_13_5_io_out_weight),
    .io_out_psum(PE_Array_13_5_io_out_psum)
  );
  basic_PE PE_Array_13_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_6_clock),
    .reset(PE_Array_13_6_reset),
    .io_in_activate(PE_Array_13_6_io_in_activate),
    .io_in_weight(PE_Array_13_6_io_in_weight),
    .io_in_psum(PE_Array_13_6_io_in_psum),
    .io_in_flow(PE_Array_13_6_io_in_flow),
    .io_in_shift(PE_Array_13_6_io_in_shift),
    .io_out_activate(PE_Array_13_6_io_out_activate),
    .io_out_weight(PE_Array_13_6_io_out_weight),
    .io_out_psum(PE_Array_13_6_io_out_psum)
  );
  basic_PE PE_Array_13_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_7_clock),
    .reset(PE_Array_13_7_reset),
    .io_in_activate(PE_Array_13_7_io_in_activate),
    .io_in_weight(PE_Array_13_7_io_in_weight),
    .io_in_psum(PE_Array_13_7_io_in_psum),
    .io_in_flow(PE_Array_13_7_io_in_flow),
    .io_in_shift(PE_Array_13_7_io_in_shift),
    .io_out_activate(PE_Array_13_7_io_out_activate),
    .io_out_weight(PE_Array_13_7_io_out_weight),
    .io_out_psum(PE_Array_13_7_io_out_psum)
  );
  basic_PE PE_Array_13_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_8_clock),
    .reset(PE_Array_13_8_reset),
    .io_in_activate(PE_Array_13_8_io_in_activate),
    .io_in_weight(PE_Array_13_8_io_in_weight),
    .io_in_psum(PE_Array_13_8_io_in_psum),
    .io_in_flow(PE_Array_13_8_io_in_flow),
    .io_in_shift(PE_Array_13_8_io_in_shift),
    .io_out_activate(PE_Array_13_8_io_out_activate),
    .io_out_weight(PE_Array_13_8_io_out_weight),
    .io_out_psum(PE_Array_13_8_io_out_psum)
  );
  basic_PE PE_Array_13_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_9_clock),
    .reset(PE_Array_13_9_reset),
    .io_in_activate(PE_Array_13_9_io_in_activate),
    .io_in_weight(PE_Array_13_9_io_in_weight),
    .io_in_psum(PE_Array_13_9_io_in_psum),
    .io_in_flow(PE_Array_13_9_io_in_flow),
    .io_in_shift(PE_Array_13_9_io_in_shift),
    .io_out_activate(PE_Array_13_9_io_out_activate),
    .io_out_weight(PE_Array_13_9_io_out_weight),
    .io_out_psum(PE_Array_13_9_io_out_psum)
  );
  basic_PE PE_Array_13_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_10_clock),
    .reset(PE_Array_13_10_reset),
    .io_in_activate(PE_Array_13_10_io_in_activate),
    .io_in_weight(PE_Array_13_10_io_in_weight),
    .io_in_psum(PE_Array_13_10_io_in_psum),
    .io_in_flow(PE_Array_13_10_io_in_flow),
    .io_in_shift(PE_Array_13_10_io_in_shift),
    .io_out_activate(PE_Array_13_10_io_out_activate),
    .io_out_weight(PE_Array_13_10_io_out_weight),
    .io_out_psum(PE_Array_13_10_io_out_psum)
  );
  basic_PE PE_Array_13_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_11_clock),
    .reset(PE_Array_13_11_reset),
    .io_in_activate(PE_Array_13_11_io_in_activate),
    .io_in_weight(PE_Array_13_11_io_in_weight),
    .io_in_psum(PE_Array_13_11_io_in_psum),
    .io_in_flow(PE_Array_13_11_io_in_flow),
    .io_in_shift(PE_Array_13_11_io_in_shift),
    .io_out_activate(PE_Array_13_11_io_out_activate),
    .io_out_weight(PE_Array_13_11_io_out_weight),
    .io_out_psum(PE_Array_13_11_io_out_psum)
  );
  basic_PE PE_Array_13_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_12_clock),
    .reset(PE_Array_13_12_reset),
    .io_in_activate(PE_Array_13_12_io_in_activate),
    .io_in_weight(PE_Array_13_12_io_in_weight),
    .io_in_psum(PE_Array_13_12_io_in_psum),
    .io_in_flow(PE_Array_13_12_io_in_flow),
    .io_in_shift(PE_Array_13_12_io_in_shift),
    .io_out_activate(PE_Array_13_12_io_out_activate),
    .io_out_weight(PE_Array_13_12_io_out_weight),
    .io_out_psum(PE_Array_13_12_io_out_psum)
  );
  basic_PE PE_Array_13_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_13_clock),
    .reset(PE_Array_13_13_reset),
    .io_in_activate(PE_Array_13_13_io_in_activate),
    .io_in_weight(PE_Array_13_13_io_in_weight),
    .io_in_psum(PE_Array_13_13_io_in_psum),
    .io_in_flow(PE_Array_13_13_io_in_flow),
    .io_in_shift(PE_Array_13_13_io_in_shift),
    .io_out_activate(PE_Array_13_13_io_out_activate),
    .io_out_weight(PE_Array_13_13_io_out_weight),
    .io_out_psum(PE_Array_13_13_io_out_psum)
  );
  basic_PE PE_Array_13_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_14_clock),
    .reset(PE_Array_13_14_reset),
    .io_in_activate(PE_Array_13_14_io_in_activate),
    .io_in_weight(PE_Array_13_14_io_in_weight),
    .io_in_psum(PE_Array_13_14_io_in_psum),
    .io_in_flow(PE_Array_13_14_io_in_flow),
    .io_in_shift(PE_Array_13_14_io_in_shift),
    .io_out_activate(PE_Array_13_14_io_out_activate),
    .io_out_weight(PE_Array_13_14_io_out_weight),
    .io_out_psum(PE_Array_13_14_io_out_psum)
  );
  basic_PE PE_Array_13_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_15_clock),
    .reset(PE_Array_13_15_reset),
    .io_in_activate(PE_Array_13_15_io_in_activate),
    .io_in_weight(PE_Array_13_15_io_in_weight),
    .io_in_psum(PE_Array_13_15_io_in_psum),
    .io_in_flow(PE_Array_13_15_io_in_flow),
    .io_in_shift(PE_Array_13_15_io_in_shift),
    .io_out_activate(PE_Array_13_15_io_out_activate),
    .io_out_weight(PE_Array_13_15_io_out_weight),
    .io_out_psum(PE_Array_13_15_io_out_psum)
  );
  basic_PE PE_Array_14_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_0_clock),
    .reset(PE_Array_14_0_reset),
    .io_in_activate(PE_Array_14_0_io_in_activate),
    .io_in_weight(PE_Array_14_0_io_in_weight),
    .io_in_psum(PE_Array_14_0_io_in_psum),
    .io_in_flow(PE_Array_14_0_io_in_flow),
    .io_in_shift(PE_Array_14_0_io_in_shift),
    .io_out_activate(PE_Array_14_0_io_out_activate),
    .io_out_weight(PE_Array_14_0_io_out_weight),
    .io_out_psum(PE_Array_14_0_io_out_psum)
  );
  basic_PE PE_Array_14_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_1_clock),
    .reset(PE_Array_14_1_reset),
    .io_in_activate(PE_Array_14_1_io_in_activate),
    .io_in_weight(PE_Array_14_1_io_in_weight),
    .io_in_psum(PE_Array_14_1_io_in_psum),
    .io_in_flow(PE_Array_14_1_io_in_flow),
    .io_in_shift(PE_Array_14_1_io_in_shift),
    .io_out_activate(PE_Array_14_1_io_out_activate),
    .io_out_weight(PE_Array_14_1_io_out_weight),
    .io_out_psum(PE_Array_14_1_io_out_psum)
  );
  basic_PE PE_Array_14_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_2_clock),
    .reset(PE_Array_14_2_reset),
    .io_in_activate(PE_Array_14_2_io_in_activate),
    .io_in_weight(PE_Array_14_2_io_in_weight),
    .io_in_psum(PE_Array_14_2_io_in_psum),
    .io_in_flow(PE_Array_14_2_io_in_flow),
    .io_in_shift(PE_Array_14_2_io_in_shift),
    .io_out_activate(PE_Array_14_2_io_out_activate),
    .io_out_weight(PE_Array_14_2_io_out_weight),
    .io_out_psum(PE_Array_14_2_io_out_psum)
  );
  basic_PE PE_Array_14_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_3_clock),
    .reset(PE_Array_14_3_reset),
    .io_in_activate(PE_Array_14_3_io_in_activate),
    .io_in_weight(PE_Array_14_3_io_in_weight),
    .io_in_psum(PE_Array_14_3_io_in_psum),
    .io_in_flow(PE_Array_14_3_io_in_flow),
    .io_in_shift(PE_Array_14_3_io_in_shift),
    .io_out_activate(PE_Array_14_3_io_out_activate),
    .io_out_weight(PE_Array_14_3_io_out_weight),
    .io_out_psum(PE_Array_14_3_io_out_psum)
  );
  basic_PE PE_Array_14_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_4_clock),
    .reset(PE_Array_14_4_reset),
    .io_in_activate(PE_Array_14_4_io_in_activate),
    .io_in_weight(PE_Array_14_4_io_in_weight),
    .io_in_psum(PE_Array_14_4_io_in_psum),
    .io_in_flow(PE_Array_14_4_io_in_flow),
    .io_in_shift(PE_Array_14_4_io_in_shift),
    .io_out_activate(PE_Array_14_4_io_out_activate),
    .io_out_weight(PE_Array_14_4_io_out_weight),
    .io_out_psum(PE_Array_14_4_io_out_psum)
  );
  basic_PE PE_Array_14_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_5_clock),
    .reset(PE_Array_14_5_reset),
    .io_in_activate(PE_Array_14_5_io_in_activate),
    .io_in_weight(PE_Array_14_5_io_in_weight),
    .io_in_psum(PE_Array_14_5_io_in_psum),
    .io_in_flow(PE_Array_14_5_io_in_flow),
    .io_in_shift(PE_Array_14_5_io_in_shift),
    .io_out_activate(PE_Array_14_5_io_out_activate),
    .io_out_weight(PE_Array_14_5_io_out_weight),
    .io_out_psum(PE_Array_14_5_io_out_psum)
  );
  basic_PE PE_Array_14_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_6_clock),
    .reset(PE_Array_14_6_reset),
    .io_in_activate(PE_Array_14_6_io_in_activate),
    .io_in_weight(PE_Array_14_6_io_in_weight),
    .io_in_psum(PE_Array_14_6_io_in_psum),
    .io_in_flow(PE_Array_14_6_io_in_flow),
    .io_in_shift(PE_Array_14_6_io_in_shift),
    .io_out_activate(PE_Array_14_6_io_out_activate),
    .io_out_weight(PE_Array_14_6_io_out_weight),
    .io_out_psum(PE_Array_14_6_io_out_psum)
  );
  basic_PE PE_Array_14_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_7_clock),
    .reset(PE_Array_14_7_reset),
    .io_in_activate(PE_Array_14_7_io_in_activate),
    .io_in_weight(PE_Array_14_7_io_in_weight),
    .io_in_psum(PE_Array_14_7_io_in_psum),
    .io_in_flow(PE_Array_14_7_io_in_flow),
    .io_in_shift(PE_Array_14_7_io_in_shift),
    .io_out_activate(PE_Array_14_7_io_out_activate),
    .io_out_weight(PE_Array_14_7_io_out_weight),
    .io_out_psum(PE_Array_14_7_io_out_psum)
  );
  basic_PE PE_Array_14_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_8_clock),
    .reset(PE_Array_14_8_reset),
    .io_in_activate(PE_Array_14_8_io_in_activate),
    .io_in_weight(PE_Array_14_8_io_in_weight),
    .io_in_psum(PE_Array_14_8_io_in_psum),
    .io_in_flow(PE_Array_14_8_io_in_flow),
    .io_in_shift(PE_Array_14_8_io_in_shift),
    .io_out_activate(PE_Array_14_8_io_out_activate),
    .io_out_weight(PE_Array_14_8_io_out_weight),
    .io_out_psum(PE_Array_14_8_io_out_psum)
  );
  basic_PE PE_Array_14_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_9_clock),
    .reset(PE_Array_14_9_reset),
    .io_in_activate(PE_Array_14_9_io_in_activate),
    .io_in_weight(PE_Array_14_9_io_in_weight),
    .io_in_psum(PE_Array_14_9_io_in_psum),
    .io_in_flow(PE_Array_14_9_io_in_flow),
    .io_in_shift(PE_Array_14_9_io_in_shift),
    .io_out_activate(PE_Array_14_9_io_out_activate),
    .io_out_weight(PE_Array_14_9_io_out_weight),
    .io_out_psum(PE_Array_14_9_io_out_psum)
  );
  basic_PE PE_Array_14_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_10_clock),
    .reset(PE_Array_14_10_reset),
    .io_in_activate(PE_Array_14_10_io_in_activate),
    .io_in_weight(PE_Array_14_10_io_in_weight),
    .io_in_psum(PE_Array_14_10_io_in_psum),
    .io_in_flow(PE_Array_14_10_io_in_flow),
    .io_in_shift(PE_Array_14_10_io_in_shift),
    .io_out_activate(PE_Array_14_10_io_out_activate),
    .io_out_weight(PE_Array_14_10_io_out_weight),
    .io_out_psum(PE_Array_14_10_io_out_psum)
  );
  basic_PE PE_Array_14_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_11_clock),
    .reset(PE_Array_14_11_reset),
    .io_in_activate(PE_Array_14_11_io_in_activate),
    .io_in_weight(PE_Array_14_11_io_in_weight),
    .io_in_psum(PE_Array_14_11_io_in_psum),
    .io_in_flow(PE_Array_14_11_io_in_flow),
    .io_in_shift(PE_Array_14_11_io_in_shift),
    .io_out_activate(PE_Array_14_11_io_out_activate),
    .io_out_weight(PE_Array_14_11_io_out_weight),
    .io_out_psum(PE_Array_14_11_io_out_psum)
  );
  basic_PE PE_Array_14_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_12_clock),
    .reset(PE_Array_14_12_reset),
    .io_in_activate(PE_Array_14_12_io_in_activate),
    .io_in_weight(PE_Array_14_12_io_in_weight),
    .io_in_psum(PE_Array_14_12_io_in_psum),
    .io_in_flow(PE_Array_14_12_io_in_flow),
    .io_in_shift(PE_Array_14_12_io_in_shift),
    .io_out_activate(PE_Array_14_12_io_out_activate),
    .io_out_weight(PE_Array_14_12_io_out_weight),
    .io_out_psum(PE_Array_14_12_io_out_psum)
  );
  basic_PE PE_Array_14_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_13_clock),
    .reset(PE_Array_14_13_reset),
    .io_in_activate(PE_Array_14_13_io_in_activate),
    .io_in_weight(PE_Array_14_13_io_in_weight),
    .io_in_psum(PE_Array_14_13_io_in_psum),
    .io_in_flow(PE_Array_14_13_io_in_flow),
    .io_in_shift(PE_Array_14_13_io_in_shift),
    .io_out_activate(PE_Array_14_13_io_out_activate),
    .io_out_weight(PE_Array_14_13_io_out_weight),
    .io_out_psum(PE_Array_14_13_io_out_psum)
  );
  basic_PE PE_Array_14_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_14_clock),
    .reset(PE_Array_14_14_reset),
    .io_in_activate(PE_Array_14_14_io_in_activate),
    .io_in_weight(PE_Array_14_14_io_in_weight),
    .io_in_psum(PE_Array_14_14_io_in_psum),
    .io_in_flow(PE_Array_14_14_io_in_flow),
    .io_in_shift(PE_Array_14_14_io_in_shift),
    .io_out_activate(PE_Array_14_14_io_out_activate),
    .io_out_weight(PE_Array_14_14_io_out_weight),
    .io_out_psum(PE_Array_14_14_io_out_psum)
  );
  basic_PE PE_Array_14_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_15_clock),
    .reset(PE_Array_14_15_reset),
    .io_in_activate(PE_Array_14_15_io_in_activate),
    .io_in_weight(PE_Array_14_15_io_in_weight),
    .io_in_psum(PE_Array_14_15_io_in_psum),
    .io_in_flow(PE_Array_14_15_io_in_flow),
    .io_in_shift(PE_Array_14_15_io_in_shift),
    .io_out_activate(PE_Array_14_15_io_out_activate),
    .io_out_weight(PE_Array_14_15_io_out_weight),
    .io_out_psum(PE_Array_14_15_io_out_psum)
  );
  basic_PE PE_Array_15_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_0_clock),
    .reset(PE_Array_15_0_reset),
    .io_in_activate(PE_Array_15_0_io_in_activate),
    .io_in_weight(PE_Array_15_0_io_in_weight),
    .io_in_psum(PE_Array_15_0_io_in_psum),
    .io_in_flow(PE_Array_15_0_io_in_flow),
    .io_in_shift(PE_Array_15_0_io_in_shift),
    .io_out_activate(PE_Array_15_0_io_out_activate),
    .io_out_weight(PE_Array_15_0_io_out_weight),
    .io_out_psum(PE_Array_15_0_io_out_psum)
  );
  basic_PE PE_Array_15_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_1_clock),
    .reset(PE_Array_15_1_reset),
    .io_in_activate(PE_Array_15_1_io_in_activate),
    .io_in_weight(PE_Array_15_1_io_in_weight),
    .io_in_psum(PE_Array_15_1_io_in_psum),
    .io_in_flow(PE_Array_15_1_io_in_flow),
    .io_in_shift(PE_Array_15_1_io_in_shift),
    .io_out_activate(PE_Array_15_1_io_out_activate),
    .io_out_weight(PE_Array_15_1_io_out_weight),
    .io_out_psum(PE_Array_15_1_io_out_psum)
  );
  basic_PE PE_Array_15_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_2_clock),
    .reset(PE_Array_15_2_reset),
    .io_in_activate(PE_Array_15_2_io_in_activate),
    .io_in_weight(PE_Array_15_2_io_in_weight),
    .io_in_psum(PE_Array_15_2_io_in_psum),
    .io_in_flow(PE_Array_15_2_io_in_flow),
    .io_in_shift(PE_Array_15_2_io_in_shift),
    .io_out_activate(PE_Array_15_2_io_out_activate),
    .io_out_weight(PE_Array_15_2_io_out_weight),
    .io_out_psum(PE_Array_15_2_io_out_psum)
  );
  basic_PE PE_Array_15_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_3_clock),
    .reset(PE_Array_15_3_reset),
    .io_in_activate(PE_Array_15_3_io_in_activate),
    .io_in_weight(PE_Array_15_3_io_in_weight),
    .io_in_psum(PE_Array_15_3_io_in_psum),
    .io_in_flow(PE_Array_15_3_io_in_flow),
    .io_in_shift(PE_Array_15_3_io_in_shift),
    .io_out_activate(PE_Array_15_3_io_out_activate),
    .io_out_weight(PE_Array_15_3_io_out_weight),
    .io_out_psum(PE_Array_15_3_io_out_psum)
  );
  basic_PE PE_Array_15_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_4_clock),
    .reset(PE_Array_15_4_reset),
    .io_in_activate(PE_Array_15_4_io_in_activate),
    .io_in_weight(PE_Array_15_4_io_in_weight),
    .io_in_psum(PE_Array_15_4_io_in_psum),
    .io_in_flow(PE_Array_15_4_io_in_flow),
    .io_in_shift(PE_Array_15_4_io_in_shift),
    .io_out_activate(PE_Array_15_4_io_out_activate),
    .io_out_weight(PE_Array_15_4_io_out_weight),
    .io_out_psum(PE_Array_15_4_io_out_psum)
  );
  basic_PE PE_Array_15_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_5_clock),
    .reset(PE_Array_15_5_reset),
    .io_in_activate(PE_Array_15_5_io_in_activate),
    .io_in_weight(PE_Array_15_5_io_in_weight),
    .io_in_psum(PE_Array_15_5_io_in_psum),
    .io_in_flow(PE_Array_15_5_io_in_flow),
    .io_in_shift(PE_Array_15_5_io_in_shift),
    .io_out_activate(PE_Array_15_5_io_out_activate),
    .io_out_weight(PE_Array_15_5_io_out_weight),
    .io_out_psum(PE_Array_15_5_io_out_psum)
  );
  basic_PE PE_Array_15_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_6_clock),
    .reset(PE_Array_15_6_reset),
    .io_in_activate(PE_Array_15_6_io_in_activate),
    .io_in_weight(PE_Array_15_6_io_in_weight),
    .io_in_psum(PE_Array_15_6_io_in_psum),
    .io_in_flow(PE_Array_15_6_io_in_flow),
    .io_in_shift(PE_Array_15_6_io_in_shift),
    .io_out_activate(PE_Array_15_6_io_out_activate),
    .io_out_weight(PE_Array_15_6_io_out_weight),
    .io_out_psum(PE_Array_15_6_io_out_psum)
  );
  basic_PE PE_Array_15_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_7_clock),
    .reset(PE_Array_15_7_reset),
    .io_in_activate(PE_Array_15_7_io_in_activate),
    .io_in_weight(PE_Array_15_7_io_in_weight),
    .io_in_psum(PE_Array_15_7_io_in_psum),
    .io_in_flow(PE_Array_15_7_io_in_flow),
    .io_in_shift(PE_Array_15_7_io_in_shift),
    .io_out_activate(PE_Array_15_7_io_out_activate),
    .io_out_weight(PE_Array_15_7_io_out_weight),
    .io_out_psum(PE_Array_15_7_io_out_psum)
  );
  basic_PE PE_Array_15_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_8_clock),
    .reset(PE_Array_15_8_reset),
    .io_in_activate(PE_Array_15_8_io_in_activate),
    .io_in_weight(PE_Array_15_8_io_in_weight),
    .io_in_psum(PE_Array_15_8_io_in_psum),
    .io_in_flow(PE_Array_15_8_io_in_flow),
    .io_in_shift(PE_Array_15_8_io_in_shift),
    .io_out_activate(PE_Array_15_8_io_out_activate),
    .io_out_weight(PE_Array_15_8_io_out_weight),
    .io_out_psum(PE_Array_15_8_io_out_psum)
  );
  basic_PE PE_Array_15_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_9_clock),
    .reset(PE_Array_15_9_reset),
    .io_in_activate(PE_Array_15_9_io_in_activate),
    .io_in_weight(PE_Array_15_9_io_in_weight),
    .io_in_psum(PE_Array_15_9_io_in_psum),
    .io_in_flow(PE_Array_15_9_io_in_flow),
    .io_in_shift(PE_Array_15_9_io_in_shift),
    .io_out_activate(PE_Array_15_9_io_out_activate),
    .io_out_weight(PE_Array_15_9_io_out_weight),
    .io_out_psum(PE_Array_15_9_io_out_psum)
  );
  basic_PE PE_Array_15_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_10_clock),
    .reset(PE_Array_15_10_reset),
    .io_in_activate(PE_Array_15_10_io_in_activate),
    .io_in_weight(PE_Array_15_10_io_in_weight),
    .io_in_psum(PE_Array_15_10_io_in_psum),
    .io_in_flow(PE_Array_15_10_io_in_flow),
    .io_in_shift(PE_Array_15_10_io_in_shift),
    .io_out_activate(PE_Array_15_10_io_out_activate),
    .io_out_weight(PE_Array_15_10_io_out_weight),
    .io_out_psum(PE_Array_15_10_io_out_psum)
  );
  basic_PE PE_Array_15_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_11_clock),
    .reset(PE_Array_15_11_reset),
    .io_in_activate(PE_Array_15_11_io_in_activate),
    .io_in_weight(PE_Array_15_11_io_in_weight),
    .io_in_psum(PE_Array_15_11_io_in_psum),
    .io_in_flow(PE_Array_15_11_io_in_flow),
    .io_in_shift(PE_Array_15_11_io_in_shift),
    .io_out_activate(PE_Array_15_11_io_out_activate),
    .io_out_weight(PE_Array_15_11_io_out_weight),
    .io_out_psum(PE_Array_15_11_io_out_psum)
  );
  basic_PE PE_Array_15_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_12_clock),
    .reset(PE_Array_15_12_reset),
    .io_in_activate(PE_Array_15_12_io_in_activate),
    .io_in_weight(PE_Array_15_12_io_in_weight),
    .io_in_psum(PE_Array_15_12_io_in_psum),
    .io_in_flow(PE_Array_15_12_io_in_flow),
    .io_in_shift(PE_Array_15_12_io_in_shift),
    .io_out_activate(PE_Array_15_12_io_out_activate),
    .io_out_weight(PE_Array_15_12_io_out_weight),
    .io_out_psum(PE_Array_15_12_io_out_psum)
  );
  basic_PE PE_Array_15_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_13_clock),
    .reset(PE_Array_15_13_reset),
    .io_in_activate(PE_Array_15_13_io_in_activate),
    .io_in_weight(PE_Array_15_13_io_in_weight),
    .io_in_psum(PE_Array_15_13_io_in_psum),
    .io_in_flow(PE_Array_15_13_io_in_flow),
    .io_in_shift(PE_Array_15_13_io_in_shift),
    .io_out_activate(PE_Array_15_13_io_out_activate),
    .io_out_weight(PE_Array_15_13_io_out_weight),
    .io_out_psum(PE_Array_15_13_io_out_psum)
  );
  basic_PE PE_Array_15_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_14_clock),
    .reset(PE_Array_15_14_reset),
    .io_in_activate(PE_Array_15_14_io_in_activate),
    .io_in_weight(PE_Array_15_14_io_in_weight),
    .io_in_psum(PE_Array_15_14_io_in_psum),
    .io_in_flow(PE_Array_15_14_io_in_flow),
    .io_in_shift(PE_Array_15_14_io_in_shift),
    .io_out_activate(PE_Array_15_14_io_out_activate),
    .io_out_weight(PE_Array_15_14_io_out_weight),
    .io_out_psum(PE_Array_15_14_io_out_psum)
  );
  basic_PE PE_Array_15_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_15_clock),
    .reset(PE_Array_15_15_reset),
    .io_in_activate(PE_Array_15_15_io_in_activate),
    .io_in_weight(PE_Array_15_15_io_in_weight),
    .io_in_psum(PE_Array_15_15_io_in_psum),
    .io_in_flow(PE_Array_15_15_io_in_flow),
    .io_in_shift(PE_Array_15_15_io_in_shift),
    .io_out_activate(PE_Array_15_15_io_out_activate),
    .io_out_weight(PE_Array_15_15_io_out_weight),
    .io_out_psum(PE_Array_15_15_io_out_psum)
  );
  assign io_psum_0 = PE_Array_15_0_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_1 = PE_Array_15_1_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_2 = PE_Array_15_2_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_3 = PE_Array_15_3_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_4 = PE_Array_15_4_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_5 = PE_Array_15_5_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_6 = PE_Array_15_6_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_7 = PE_Array_15_7_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_8 = PE_Array_15_8_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_9 = PE_Array_15_9_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_10 = PE_Array_15_10_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_11 = PE_Array_15_11_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_12 = PE_Array_15_12_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_13 = PE_Array_15_13_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_14 = PE_Array_15_14_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_15 = PE_Array_15_15_io_out_psum; // @[DataPath.scala 24:10]
  assign io_valid_0 = valid_reg[0]; // @[Systolic_Array.scala 73:33]
  assign io_valid_1 = valid_reg[1]; // @[Systolic_Array.scala 73:33]
  assign io_valid_2 = valid_reg[2]; // @[Systolic_Array.scala 73:33]
  assign io_valid_3 = valid_reg[3]; // @[Systolic_Array.scala 73:33]
  assign io_valid_4 = valid_reg[4]; // @[Systolic_Array.scala 73:33]
  assign io_valid_5 = valid_reg[5]; // @[Systolic_Array.scala 73:33]
  assign io_valid_6 = valid_reg[6]; // @[Systolic_Array.scala 73:33]
  assign io_valid_7 = valid_reg[7]; // @[Systolic_Array.scala 73:33]
  assign io_valid_8 = valid_reg[8]; // @[Systolic_Array.scala 73:33]
  assign io_valid_9 = valid_reg[9]; // @[Systolic_Array.scala 73:33]
  assign io_valid_10 = valid_reg[10]; // @[Systolic_Array.scala 73:33]
  assign io_valid_11 = valid_reg[11]; // @[Systolic_Array.scala 73:33]
  assign io_valid_12 = valid_reg[12]; // @[Systolic_Array.scala 73:33]
  assign io_valid_13 = valid_reg[13]; // @[Systolic_Array.scala 73:33]
  assign io_valid_14 = valid_reg[14]; // @[Systolic_Array.scala 73:33]
  assign io_valid_15 = valid_reg[15]; // @[Systolic_Array.scala 73:33]
  assign PE_Array_0_0_clock = clock;
  assign PE_Array_0_0_reset = reset;
  assign PE_Array_0_0_io_in_activate = io_activate_0; // @[DataPath.scala 11:26]
  assign PE_Array_0_0_io_in_weight = io_weight_0; // @[DataPath.scala 20:23]
  assign PE_Array_0_0_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_1_clock = clock;
  assign PE_Array_0_1_reset = reset;
  assign PE_Array_0_1_io_in_activate = PE_Array_0_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_1_io_in_weight = io_weight_1; // @[DataPath.scala 20:23]
  assign PE_Array_0_1_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_2_clock = clock;
  assign PE_Array_0_2_reset = reset;
  assign PE_Array_0_2_io_in_activate = PE_Array_0_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_2_io_in_weight = io_weight_2; // @[DataPath.scala 20:23]
  assign PE_Array_0_2_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_3_clock = clock;
  assign PE_Array_0_3_reset = reset;
  assign PE_Array_0_3_io_in_activate = PE_Array_0_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_3_io_in_weight = io_weight_3; // @[DataPath.scala 20:23]
  assign PE_Array_0_3_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_4_clock = clock;
  assign PE_Array_0_4_reset = reset;
  assign PE_Array_0_4_io_in_activate = PE_Array_0_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_4_io_in_weight = io_weight_4; // @[DataPath.scala 20:23]
  assign PE_Array_0_4_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_5_clock = clock;
  assign PE_Array_0_5_reset = reset;
  assign PE_Array_0_5_io_in_activate = PE_Array_0_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_5_io_in_weight = io_weight_5; // @[DataPath.scala 20:23]
  assign PE_Array_0_5_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_6_clock = clock;
  assign PE_Array_0_6_reset = reset;
  assign PE_Array_0_6_io_in_activate = PE_Array_0_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_6_io_in_weight = io_weight_6; // @[DataPath.scala 20:23]
  assign PE_Array_0_6_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_7_clock = clock;
  assign PE_Array_0_7_reset = reset;
  assign PE_Array_0_7_io_in_activate = PE_Array_0_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_7_io_in_weight = io_weight_7; // @[DataPath.scala 20:23]
  assign PE_Array_0_7_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_8_clock = clock;
  assign PE_Array_0_8_reset = reset;
  assign PE_Array_0_8_io_in_activate = PE_Array_0_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_8_io_in_weight = io_weight_8; // @[DataPath.scala 20:23]
  assign PE_Array_0_8_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_9_clock = clock;
  assign PE_Array_0_9_reset = reset;
  assign PE_Array_0_9_io_in_activate = PE_Array_0_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_9_io_in_weight = io_weight_9; // @[DataPath.scala 20:23]
  assign PE_Array_0_9_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_10_clock = clock;
  assign PE_Array_0_10_reset = reset;
  assign PE_Array_0_10_io_in_activate = PE_Array_0_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_10_io_in_weight = io_weight_10; // @[DataPath.scala 20:23]
  assign PE_Array_0_10_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_11_clock = clock;
  assign PE_Array_0_11_reset = reset;
  assign PE_Array_0_11_io_in_activate = PE_Array_0_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_11_io_in_weight = io_weight_11; // @[DataPath.scala 20:23]
  assign PE_Array_0_11_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_12_clock = clock;
  assign PE_Array_0_12_reset = reset;
  assign PE_Array_0_12_io_in_activate = PE_Array_0_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_12_io_in_weight = io_weight_12; // @[DataPath.scala 20:23]
  assign PE_Array_0_12_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_13_clock = clock;
  assign PE_Array_0_13_reset = reset;
  assign PE_Array_0_13_io_in_activate = PE_Array_0_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_13_io_in_weight = io_weight_13; // @[DataPath.scala 20:23]
  assign PE_Array_0_13_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_14_clock = clock;
  assign PE_Array_0_14_reset = reset;
  assign PE_Array_0_14_io_in_activate = PE_Array_0_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_14_io_in_weight = io_weight_14; // @[DataPath.scala 20:23]
  assign PE_Array_0_14_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_15_clock = clock;
  assign PE_Array_0_15_reset = reset;
  assign PE_Array_0_15_io_in_activate = PE_Array_0_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_15_io_in_weight = io_weight_15; // @[DataPath.scala 20:23]
  assign PE_Array_0_15_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_0_clock = clock;
  assign PE_Array_1_0_reset = reset;
  assign PE_Array_1_0_io_in_activate = io_activate_1; // @[DataPath.scala 11:26]
  assign PE_Array_1_0_io_in_weight = PE_Array_0_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_0_io_in_psum = PE_Array_0_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_1_clock = clock;
  assign PE_Array_1_1_reset = reset;
  assign PE_Array_1_1_io_in_activate = PE_Array_1_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_1_io_in_weight = PE_Array_0_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_1_io_in_psum = PE_Array_0_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_2_clock = clock;
  assign PE_Array_1_2_reset = reset;
  assign PE_Array_1_2_io_in_activate = PE_Array_1_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_2_io_in_weight = PE_Array_0_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_2_io_in_psum = PE_Array_0_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_3_clock = clock;
  assign PE_Array_1_3_reset = reset;
  assign PE_Array_1_3_io_in_activate = PE_Array_1_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_3_io_in_weight = PE_Array_0_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_3_io_in_psum = PE_Array_0_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_4_clock = clock;
  assign PE_Array_1_4_reset = reset;
  assign PE_Array_1_4_io_in_activate = PE_Array_1_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_4_io_in_weight = PE_Array_0_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_4_io_in_psum = PE_Array_0_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_5_clock = clock;
  assign PE_Array_1_5_reset = reset;
  assign PE_Array_1_5_io_in_activate = PE_Array_1_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_5_io_in_weight = PE_Array_0_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_5_io_in_psum = PE_Array_0_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_6_clock = clock;
  assign PE_Array_1_6_reset = reset;
  assign PE_Array_1_6_io_in_activate = PE_Array_1_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_6_io_in_weight = PE_Array_0_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_6_io_in_psum = PE_Array_0_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_7_clock = clock;
  assign PE_Array_1_7_reset = reset;
  assign PE_Array_1_7_io_in_activate = PE_Array_1_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_7_io_in_weight = PE_Array_0_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_7_io_in_psum = PE_Array_0_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_8_clock = clock;
  assign PE_Array_1_8_reset = reset;
  assign PE_Array_1_8_io_in_activate = PE_Array_1_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_8_io_in_weight = PE_Array_0_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_8_io_in_psum = PE_Array_0_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_9_clock = clock;
  assign PE_Array_1_9_reset = reset;
  assign PE_Array_1_9_io_in_activate = PE_Array_1_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_9_io_in_weight = PE_Array_0_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_9_io_in_psum = PE_Array_0_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_10_clock = clock;
  assign PE_Array_1_10_reset = reset;
  assign PE_Array_1_10_io_in_activate = PE_Array_1_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_10_io_in_weight = PE_Array_0_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_10_io_in_psum = PE_Array_0_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_11_clock = clock;
  assign PE_Array_1_11_reset = reset;
  assign PE_Array_1_11_io_in_activate = PE_Array_1_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_11_io_in_weight = PE_Array_0_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_11_io_in_psum = PE_Array_0_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_12_clock = clock;
  assign PE_Array_1_12_reset = reset;
  assign PE_Array_1_12_io_in_activate = PE_Array_1_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_12_io_in_weight = PE_Array_0_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_12_io_in_psum = PE_Array_0_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_13_clock = clock;
  assign PE_Array_1_13_reset = reset;
  assign PE_Array_1_13_io_in_activate = PE_Array_1_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_13_io_in_weight = PE_Array_0_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_13_io_in_psum = PE_Array_0_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_14_clock = clock;
  assign PE_Array_1_14_reset = reset;
  assign PE_Array_1_14_io_in_activate = PE_Array_1_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_14_io_in_weight = PE_Array_0_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_14_io_in_psum = PE_Array_0_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_15_clock = clock;
  assign PE_Array_1_15_reset = reset;
  assign PE_Array_1_15_io_in_activate = PE_Array_1_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_15_io_in_weight = PE_Array_0_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_15_io_in_psum = PE_Array_0_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_0_clock = clock;
  assign PE_Array_2_0_reset = reset;
  assign PE_Array_2_0_io_in_activate = io_activate_2; // @[DataPath.scala 11:26]
  assign PE_Array_2_0_io_in_weight = PE_Array_1_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_0_io_in_psum = PE_Array_1_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_1_clock = clock;
  assign PE_Array_2_1_reset = reset;
  assign PE_Array_2_1_io_in_activate = PE_Array_2_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_1_io_in_weight = PE_Array_1_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_1_io_in_psum = PE_Array_1_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_2_clock = clock;
  assign PE_Array_2_2_reset = reset;
  assign PE_Array_2_2_io_in_activate = PE_Array_2_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_2_io_in_weight = PE_Array_1_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_2_io_in_psum = PE_Array_1_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_3_clock = clock;
  assign PE_Array_2_3_reset = reset;
  assign PE_Array_2_3_io_in_activate = PE_Array_2_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_3_io_in_weight = PE_Array_1_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_3_io_in_psum = PE_Array_1_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_4_clock = clock;
  assign PE_Array_2_4_reset = reset;
  assign PE_Array_2_4_io_in_activate = PE_Array_2_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_4_io_in_weight = PE_Array_1_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_4_io_in_psum = PE_Array_1_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_5_clock = clock;
  assign PE_Array_2_5_reset = reset;
  assign PE_Array_2_5_io_in_activate = PE_Array_2_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_5_io_in_weight = PE_Array_1_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_5_io_in_psum = PE_Array_1_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_6_clock = clock;
  assign PE_Array_2_6_reset = reset;
  assign PE_Array_2_6_io_in_activate = PE_Array_2_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_6_io_in_weight = PE_Array_1_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_6_io_in_psum = PE_Array_1_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_7_clock = clock;
  assign PE_Array_2_7_reset = reset;
  assign PE_Array_2_7_io_in_activate = PE_Array_2_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_7_io_in_weight = PE_Array_1_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_7_io_in_psum = PE_Array_1_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_8_clock = clock;
  assign PE_Array_2_8_reset = reset;
  assign PE_Array_2_8_io_in_activate = PE_Array_2_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_8_io_in_weight = PE_Array_1_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_8_io_in_psum = PE_Array_1_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_9_clock = clock;
  assign PE_Array_2_9_reset = reset;
  assign PE_Array_2_9_io_in_activate = PE_Array_2_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_9_io_in_weight = PE_Array_1_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_9_io_in_psum = PE_Array_1_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_10_clock = clock;
  assign PE_Array_2_10_reset = reset;
  assign PE_Array_2_10_io_in_activate = PE_Array_2_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_10_io_in_weight = PE_Array_1_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_10_io_in_psum = PE_Array_1_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_11_clock = clock;
  assign PE_Array_2_11_reset = reset;
  assign PE_Array_2_11_io_in_activate = PE_Array_2_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_11_io_in_weight = PE_Array_1_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_11_io_in_psum = PE_Array_1_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_12_clock = clock;
  assign PE_Array_2_12_reset = reset;
  assign PE_Array_2_12_io_in_activate = PE_Array_2_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_12_io_in_weight = PE_Array_1_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_12_io_in_psum = PE_Array_1_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_13_clock = clock;
  assign PE_Array_2_13_reset = reset;
  assign PE_Array_2_13_io_in_activate = PE_Array_2_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_13_io_in_weight = PE_Array_1_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_13_io_in_psum = PE_Array_1_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_14_clock = clock;
  assign PE_Array_2_14_reset = reset;
  assign PE_Array_2_14_io_in_activate = PE_Array_2_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_14_io_in_weight = PE_Array_1_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_14_io_in_psum = PE_Array_1_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_15_clock = clock;
  assign PE_Array_2_15_reset = reset;
  assign PE_Array_2_15_io_in_activate = PE_Array_2_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_15_io_in_weight = PE_Array_1_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_15_io_in_psum = PE_Array_1_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_0_clock = clock;
  assign PE_Array_3_0_reset = reset;
  assign PE_Array_3_0_io_in_activate = io_activate_3; // @[DataPath.scala 11:26]
  assign PE_Array_3_0_io_in_weight = PE_Array_2_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_0_io_in_psum = PE_Array_2_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_1_clock = clock;
  assign PE_Array_3_1_reset = reset;
  assign PE_Array_3_1_io_in_activate = PE_Array_3_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_1_io_in_weight = PE_Array_2_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_1_io_in_psum = PE_Array_2_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_2_clock = clock;
  assign PE_Array_3_2_reset = reset;
  assign PE_Array_3_2_io_in_activate = PE_Array_3_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_2_io_in_weight = PE_Array_2_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_2_io_in_psum = PE_Array_2_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_3_clock = clock;
  assign PE_Array_3_3_reset = reset;
  assign PE_Array_3_3_io_in_activate = PE_Array_3_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_3_io_in_weight = PE_Array_2_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_3_io_in_psum = PE_Array_2_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_4_clock = clock;
  assign PE_Array_3_4_reset = reset;
  assign PE_Array_3_4_io_in_activate = PE_Array_3_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_4_io_in_weight = PE_Array_2_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_4_io_in_psum = PE_Array_2_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_5_clock = clock;
  assign PE_Array_3_5_reset = reset;
  assign PE_Array_3_5_io_in_activate = PE_Array_3_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_5_io_in_weight = PE_Array_2_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_5_io_in_psum = PE_Array_2_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_6_clock = clock;
  assign PE_Array_3_6_reset = reset;
  assign PE_Array_3_6_io_in_activate = PE_Array_3_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_6_io_in_weight = PE_Array_2_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_6_io_in_psum = PE_Array_2_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_7_clock = clock;
  assign PE_Array_3_7_reset = reset;
  assign PE_Array_3_7_io_in_activate = PE_Array_3_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_7_io_in_weight = PE_Array_2_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_7_io_in_psum = PE_Array_2_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_8_clock = clock;
  assign PE_Array_3_8_reset = reset;
  assign PE_Array_3_8_io_in_activate = PE_Array_3_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_8_io_in_weight = PE_Array_2_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_8_io_in_psum = PE_Array_2_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_9_clock = clock;
  assign PE_Array_3_9_reset = reset;
  assign PE_Array_3_9_io_in_activate = PE_Array_3_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_9_io_in_weight = PE_Array_2_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_9_io_in_psum = PE_Array_2_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_10_clock = clock;
  assign PE_Array_3_10_reset = reset;
  assign PE_Array_3_10_io_in_activate = PE_Array_3_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_10_io_in_weight = PE_Array_2_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_10_io_in_psum = PE_Array_2_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_11_clock = clock;
  assign PE_Array_3_11_reset = reset;
  assign PE_Array_3_11_io_in_activate = PE_Array_3_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_11_io_in_weight = PE_Array_2_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_11_io_in_psum = PE_Array_2_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_12_clock = clock;
  assign PE_Array_3_12_reset = reset;
  assign PE_Array_3_12_io_in_activate = PE_Array_3_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_12_io_in_weight = PE_Array_2_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_12_io_in_psum = PE_Array_2_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_13_clock = clock;
  assign PE_Array_3_13_reset = reset;
  assign PE_Array_3_13_io_in_activate = PE_Array_3_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_13_io_in_weight = PE_Array_2_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_13_io_in_psum = PE_Array_2_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_14_clock = clock;
  assign PE_Array_3_14_reset = reset;
  assign PE_Array_3_14_io_in_activate = PE_Array_3_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_14_io_in_weight = PE_Array_2_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_14_io_in_psum = PE_Array_2_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_15_clock = clock;
  assign PE_Array_3_15_reset = reset;
  assign PE_Array_3_15_io_in_activate = PE_Array_3_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_15_io_in_weight = PE_Array_2_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_15_io_in_psum = PE_Array_2_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_0_clock = clock;
  assign PE_Array_4_0_reset = reset;
  assign PE_Array_4_0_io_in_activate = io_activate_4; // @[DataPath.scala 11:26]
  assign PE_Array_4_0_io_in_weight = PE_Array_3_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_0_io_in_psum = PE_Array_3_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_1_clock = clock;
  assign PE_Array_4_1_reset = reset;
  assign PE_Array_4_1_io_in_activate = PE_Array_4_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_1_io_in_weight = PE_Array_3_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_1_io_in_psum = PE_Array_3_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_2_clock = clock;
  assign PE_Array_4_2_reset = reset;
  assign PE_Array_4_2_io_in_activate = PE_Array_4_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_2_io_in_weight = PE_Array_3_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_2_io_in_psum = PE_Array_3_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_3_clock = clock;
  assign PE_Array_4_3_reset = reset;
  assign PE_Array_4_3_io_in_activate = PE_Array_4_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_3_io_in_weight = PE_Array_3_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_3_io_in_psum = PE_Array_3_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_4_clock = clock;
  assign PE_Array_4_4_reset = reset;
  assign PE_Array_4_4_io_in_activate = PE_Array_4_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_4_io_in_weight = PE_Array_3_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_4_io_in_psum = PE_Array_3_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_5_clock = clock;
  assign PE_Array_4_5_reset = reset;
  assign PE_Array_4_5_io_in_activate = PE_Array_4_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_5_io_in_weight = PE_Array_3_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_5_io_in_psum = PE_Array_3_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_6_clock = clock;
  assign PE_Array_4_6_reset = reset;
  assign PE_Array_4_6_io_in_activate = PE_Array_4_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_6_io_in_weight = PE_Array_3_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_6_io_in_psum = PE_Array_3_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_7_clock = clock;
  assign PE_Array_4_7_reset = reset;
  assign PE_Array_4_7_io_in_activate = PE_Array_4_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_7_io_in_weight = PE_Array_3_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_7_io_in_psum = PE_Array_3_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_8_clock = clock;
  assign PE_Array_4_8_reset = reset;
  assign PE_Array_4_8_io_in_activate = PE_Array_4_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_8_io_in_weight = PE_Array_3_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_8_io_in_psum = PE_Array_3_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_9_clock = clock;
  assign PE_Array_4_9_reset = reset;
  assign PE_Array_4_9_io_in_activate = PE_Array_4_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_9_io_in_weight = PE_Array_3_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_9_io_in_psum = PE_Array_3_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_10_clock = clock;
  assign PE_Array_4_10_reset = reset;
  assign PE_Array_4_10_io_in_activate = PE_Array_4_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_10_io_in_weight = PE_Array_3_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_10_io_in_psum = PE_Array_3_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_11_clock = clock;
  assign PE_Array_4_11_reset = reset;
  assign PE_Array_4_11_io_in_activate = PE_Array_4_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_11_io_in_weight = PE_Array_3_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_11_io_in_psum = PE_Array_3_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_12_clock = clock;
  assign PE_Array_4_12_reset = reset;
  assign PE_Array_4_12_io_in_activate = PE_Array_4_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_12_io_in_weight = PE_Array_3_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_12_io_in_psum = PE_Array_3_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_13_clock = clock;
  assign PE_Array_4_13_reset = reset;
  assign PE_Array_4_13_io_in_activate = PE_Array_4_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_13_io_in_weight = PE_Array_3_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_13_io_in_psum = PE_Array_3_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_14_clock = clock;
  assign PE_Array_4_14_reset = reset;
  assign PE_Array_4_14_io_in_activate = PE_Array_4_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_14_io_in_weight = PE_Array_3_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_14_io_in_psum = PE_Array_3_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_15_clock = clock;
  assign PE_Array_4_15_reset = reset;
  assign PE_Array_4_15_io_in_activate = PE_Array_4_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_15_io_in_weight = PE_Array_3_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_15_io_in_psum = PE_Array_3_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_0_clock = clock;
  assign PE_Array_5_0_reset = reset;
  assign PE_Array_5_0_io_in_activate = io_activate_5; // @[DataPath.scala 11:26]
  assign PE_Array_5_0_io_in_weight = PE_Array_4_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_0_io_in_psum = PE_Array_4_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_1_clock = clock;
  assign PE_Array_5_1_reset = reset;
  assign PE_Array_5_1_io_in_activate = PE_Array_5_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_1_io_in_weight = PE_Array_4_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_1_io_in_psum = PE_Array_4_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_2_clock = clock;
  assign PE_Array_5_2_reset = reset;
  assign PE_Array_5_2_io_in_activate = PE_Array_5_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_2_io_in_weight = PE_Array_4_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_2_io_in_psum = PE_Array_4_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_3_clock = clock;
  assign PE_Array_5_3_reset = reset;
  assign PE_Array_5_3_io_in_activate = PE_Array_5_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_3_io_in_weight = PE_Array_4_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_3_io_in_psum = PE_Array_4_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_4_clock = clock;
  assign PE_Array_5_4_reset = reset;
  assign PE_Array_5_4_io_in_activate = PE_Array_5_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_4_io_in_weight = PE_Array_4_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_4_io_in_psum = PE_Array_4_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_5_clock = clock;
  assign PE_Array_5_5_reset = reset;
  assign PE_Array_5_5_io_in_activate = PE_Array_5_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_5_io_in_weight = PE_Array_4_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_5_io_in_psum = PE_Array_4_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_6_clock = clock;
  assign PE_Array_5_6_reset = reset;
  assign PE_Array_5_6_io_in_activate = PE_Array_5_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_6_io_in_weight = PE_Array_4_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_6_io_in_psum = PE_Array_4_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_7_clock = clock;
  assign PE_Array_5_7_reset = reset;
  assign PE_Array_5_7_io_in_activate = PE_Array_5_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_7_io_in_weight = PE_Array_4_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_7_io_in_psum = PE_Array_4_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_8_clock = clock;
  assign PE_Array_5_8_reset = reset;
  assign PE_Array_5_8_io_in_activate = PE_Array_5_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_8_io_in_weight = PE_Array_4_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_8_io_in_psum = PE_Array_4_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_9_clock = clock;
  assign PE_Array_5_9_reset = reset;
  assign PE_Array_5_9_io_in_activate = PE_Array_5_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_9_io_in_weight = PE_Array_4_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_9_io_in_psum = PE_Array_4_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_10_clock = clock;
  assign PE_Array_5_10_reset = reset;
  assign PE_Array_5_10_io_in_activate = PE_Array_5_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_10_io_in_weight = PE_Array_4_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_10_io_in_psum = PE_Array_4_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_11_clock = clock;
  assign PE_Array_5_11_reset = reset;
  assign PE_Array_5_11_io_in_activate = PE_Array_5_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_11_io_in_weight = PE_Array_4_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_11_io_in_psum = PE_Array_4_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_12_clock = clock;
  assign PE_Array_5_12_reset = reset;
  assign PE_Array_5_12_io_in_activate = PE_Array_5_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_12_io_in_weight = PE_Array_4_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_12_io_in_psum = PE_Array_4_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_13_clock = clock;
  assign PE_Array_5_13_reset = reset;
  assign PE_Array_5_13_io_in_activate = PE_Array_5_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_13_io_in_weight = PE_Array_4_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_13_io_in_psum = PE_Array_4_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_14_clock = clock;
  assign PE_Array_5_14_reset = reset;
  assign PE_Array_5_14_io_in_activate = PE_Array_5_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_14_io_in_weight = PE_Array_4_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_14_io_in_psum = PE_Array_4_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_15_clock = clock;
  assign PE_Array_5_15_reset = reset;
  assign PE_Array_5_15_io_in_activate = PE_Array_5_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_15_io_in_weight = PE_Array_4_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_15_io_in_psum = PE_Array_4_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_0_clock = clock;
  assign PE_Array_6_0_reset = reset;
  assign PE_Array_6_0_io_in_activate = io_activate_6; // @[DataPath.scala 11:26]
  assign PE_Array_6_0_io_in_weight = PE_Array_5_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_0_io_in_psum = PE_Array_5_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_1_clock = clock;
  assign PE_Array_6_1_reset = reset;
  assign PE_Array_6_1_io_in_activate = PE_Array_6_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_1_io_in_weight = PE_Array_5_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_1_io_in_psum = PE_Array_5_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_2_clock = clock;
  assign PE_Array_6_2_reset = reset;
  assign PE_Array_6_2_io_in_activate = PE_Array_6_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_2_io_in_weight = PE_Array_5_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_2_io_in_psum = PE_Array_5_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_3_clock = clock;
  assign PE_Array_6_3_reset = reset;
  assign PE_Array_6_3_io_in_activate = PE_Array_6_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_3_io_in_weight = PE_Array_5_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_3_io_in_psum = PE_Array_5_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_4_clock = clock;
  assign PE_Array_6_4_reset = reset;
  assign PE_Array_6_4_io_in_activate = PE_Array_6_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_4_io_in_weight = PE_Array_5_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_4_io_in_psum = PE_Array_5_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_5_clock = clock;
  assign PE_Array_6_5_reset = reset;
  assign PE_Array_6_5_io_in_activate = PE_Array_6_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_5_io_in_weight = PE_Array_5_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_5_io_in_psum = PE_Array_5_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_6_clock = clock;
  assign PE_Array_6_6_reset = reset;
  assign PE_Array_6_6_io_in_activate = PE_Array_6_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_6_io_in_weight = PE_Array_5_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_6_io_in_psum = PE_Array_5_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_7_clock = clock;
  assign PE_Array_6_7_reset = reset;
  assign PE_Array_6_7_io_in_activate = PE_Array_6_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_7_io_in_weight = PE_Array_5_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_7_io_in_psum = PE_Array_5_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_8_clock = clock;
  assign PE_Array_6_8_reset = reset;
  assign PE_Array_6_8_io_in_activate = PE_Array_6_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_8_io_in_weight = PE_Array_5_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_8_io_in_psum = PE_Array_5_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_9_clock = clock;
  assign PE_Array_6_9_reset = reset;
  assign PE_Array_6_9_io_in_activate = PE_Array_6_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_9_io_in_weight = PE_Array_5_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_9_io_in_psum = PE_Array_5_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_10_clock = clock;
  assign PE_Array_6_10_reset = reset;
  assign PE_Array_6_10_io_in_activate = PE_Array_6_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_10_io_in_weight = PE_Array_5_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_10_io_in_psum = PE_Array_5_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_11_clock = clock;
  assign PE_Array_6_11_reset = reset;
  assign PE_Array_6_11_io_in_activate = PE_Array_6_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_11_io_in_weight = PE_Array_5_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_11_io_in_psum = PE_Array_5_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_12_clock = clock;
  assign PE_Array_6_12_reset = reset;
  assign PE_Array_6_12_io_in_activate = PE_Array_6_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_12_io_in_weight = PE_Array_5_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_12_io_in_psum = PE_Array_5_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_13_clock = clock;
  assign PE_Array_6_13_reset = reset;
  assign PE_Array_6_13_io_in_activate = PE_Array_6_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_13_io_in_weight = PE_Array_5_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_13_io_in_psum = PE_Array_5_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_14_clock = clock;
  assign PE_Array_6_14_reset = reset;
  assign PE_Array_6_14_io_in_activate = PE_Array_6_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_14_io_in_weight = PE_Array_5_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_14_io_in_psum = PE_Array_5_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_15_clock = clock;
  assign PE_Array_6_15_reset = reset;
  assign PE_Array_6_15_io_in_activate = PE_Array_6_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_15_io_in_weight = PE_Array_5_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_15_io_in_psum = PE_Array_5_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_0_clock = clock;
  assign PE_Array_7_0_reset = reset;
  assign PE_Array_7_0_io_in_activate = io_activate_7; // @[DataPath.scala 11:26]
  assign PE_Array_7_0_io_in_weight = PE_Array_6_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_0_io_in_psum = PE_Array_6_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_1_clock = clock;
  assign PE_Array_7_1_reset = reset;
  assign PE_Array_7_1_io_in_activate = PE_Array_7_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_1_io_in_weight = PE_Array_6_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_1_io_in_psum = PE_Array_6_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_2_clock = clock;
  assign PE_Array_7_2_reset = reset;
  assign PE_Array_7_2_io_in_activate = PE_Array_7_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_2_io_in_weight = PE_Array_6_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_2_io_in_psum = PE_Array_6_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_3_clock = clock;
  assign PE_Array_7_3_reset = reset;
  assign PE_Array_7_3_io_in_activate = PE_Array_7_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_3_io_in_weight = PE_Array_6_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_3_io_in_psum = PE_Array_6_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_4_clock = clock;
  assign PE_Array_7_4_reset = reset;
  assign PE_Array_7_4_io_in_activate = PE_Array_7_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_4_io_in_weight = PE_Array_6_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_4_io_in_psum = PE_Array_6_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_5_clock = clock;
  assign PE_Array_7_5_reset = reset;
  assign PE_Array_7_5_io_in_activate = PE_Array_7_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_5_io_in_weight = PE_Array_6_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_5_io_in_psum = PE_Array_6_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_6_clock = clock;
  assign PE_Array_7_6_reset = reset;
  assign PE_Array_7_6_io_in_activate = PE_Array_7_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_6_io_in_weight = PE_Array_6_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_6_io_in_psum = PE_Array_6_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_7_clock = clock;
  assign PE_Array_7_7_reset = reset;
  assign PE_Array_7_7_io_in_activate = PE_Array_7_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_7_io_in_weight = PE_Array_6_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_7_io_in_psum = PE_Array_6_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_8_clock = clock;
  assign PE_Array_7_8_reset = reset;
  assign PE_Array_7_8_io_in_activate = PE_Array_7_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_8_io_in_weight = PE_Array_6_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_8_io_in_psum = PE_Array_6_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_9_clock = clock;
  assign PE_Array_7_9_reset = reset;
  assign PE_Array_7_9_io_in_activate = PE_Array_7_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_9_io_in_weight = PE_Array_6_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_9_io_in_psum = PE_Array_6_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_10_clock = clock;
  assign PE_Array_7_10_reset = reset;
  assign PE_Array_7_10_io_in_activate = PE_Array_7_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_10_io_in_weight = PE_Array_6_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_10_io_in_psum = PE_Array_6_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_11_clock = clock;
  assign PE_Array_7_11_reset = reset;
  assign PE_Array_7_11_io_in_activate = PE_Array_7_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_11_io_in_weight = PE_Array_6_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_11_io_in_psum = PE_Array_6_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_12_clock = clock;
  assign PE_Array_7_12_reset = reset;
  assign PE_Array_7_12_io_in_activate = PE_Array_7_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_12_io_in_weight = PE_Array_6_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_12_io_in_psum = PE_Array_6_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_13_clock = clock;
  assign PE_Array_7_13_reset = reset;
  assign PE_Array_7_13_io_in_activate = PE_Array_7_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_13_io_in_weight = PE_Array_6_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_13_io_in_psum = PE_Array_6_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_14_clock = clock;
  assign PE_Array_7_14_reset = reset;
  assign PE_Array_7_14_io_in_activate = PE_Array_7_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_14_io_in_weight = PE_Array_6_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_14_io_in_psum = PE_Array_6_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_15_clock = clock;
  assign PE_Array_7_15_reset = reset;
  assign PE_Array_7_15_io_in_activate = PE_Array_7_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_15_io_in_weight = PE_Array_6_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_15_io_in_psum = PE_Array_6_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_0_clock = clock;
  assign PE_Array_8_0_reset = reset;
  assign PE_Array_8_0_io_in_activate = io_activate_8; // @[DataPath.scala 11:26]
  assign PE_Array_8_0_io_in_weight = PE_Array_7_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_0_io_in_psum = PE_Array_7_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_1_clock = clock;
  assign PE_Array_8_1_reset = reset;
  assign PE_Array_8_1_io_in_activate = PE_Array_8_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_1_io_in_weight = PE_Array_7_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_1_io_in_psum = PE_Array_7_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_2_clock = clock;
  assign PE_Array_8_2_reset = reset;
  assign PE_Array_8_2_io_in_activate = PE_Array_8_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_2_io_in_weight = PE_Array_7_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_2_io_in_psum = PE_Array_7_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_3_clock = clock;
  assign PE_Array_8_3_reset = reset;
  assign PE_Array_8_3_io_in_activate = PE_Array_8_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_3_io_in_weight = PE_Array_7_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_3_io_in_psum = PE_Array_7_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_4_clock = clock;
  assign PE_Array_8_4_reset = reset;
  assign PE_Array_8_4_io_in_activate = PE_Array_8_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_4_io_in_weight = PE_Array_7_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_4_io_in_psum = PE_Array_7_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_5_clock = clock;
  assign PE_Array_8_5_reset = reset;
  assign PE_Array_8_5_io_in_activate = PE_Array_8_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_5_io_in_weight = PE_Array_7_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_5_io_in_psum = PE_Array_7_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_6_clock = clock;
  assign PE_Array_8_6_reset = reset;
  assign PE_Array_8_6_io_in_activate = PE_Array_8_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_6_io_in_weight = PE_Array_7_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_6_io_in_psum = PE_Array_7_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_7_clock = clock;
  assign PE_Array_8_7_reset = reset;
  assign PE_Array_8_7_io_in_activate = PE_Array_8_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_7_io_in_weight = PE_Array_7_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_7_io_in_psum = PE_Array_7_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_8_clock = clock;
  assign PE_Array_8_8_reset = reset;
  assign PE_Array_8_8_io_in_activate = PE_Array_8_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_8_io_in_weight = PE_Array_7_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_8_io_in_psum = PE_Array_7_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_9_clock = clock;
  assign PE_Array_8_9_reset = reset;
  assign PE_Array_8_9_io_in_activate = PE_Array_8_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_9_io_in_weight = PE_Array_7_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_9_io_in_psum = PE_Array_7_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_10_clock = clock;
  assign PE_Array_8_10_reset = reset;
  assign PE_Array_8_10_io_in_activate = PE_Array_8_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_10_io_in_weight = PE_Array_7_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_10_io_in_psum = PE_Array_7_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_11_clock = clock;
  assign PE_Array_8_11_reset = reset;
  assign PE_Array_8_11_io_in_activate = PE_Array_8_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_11_io_in_weight = PE_Array_7_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_11_io_in_psum = PE_Array_7_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_12_clock = clock;
  assign PE_Array_8_12_reset = reset;
  assign PE_Array_8_12_io_in_activate = PE_Array_8_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_12_io_in_weight = PE_Array_7_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_12_io_in_psum = PE_Array_7_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_13_clock = clock;
  assign PE_Array_8_13_reset = reset;
  assign PE_Array_8_13_io_in_activate = PE_Array_8_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_13_io_in_weight = PE_Array_7_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_13_io_in_psum = PE_Array_7_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_14_clock = clock;
  assign PE_Array_8_14_reset = reset;
  assign PE_Array_8_14_io_in_activate = PE_Array_8_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_14_io_in_weight = PE_Array_7_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_14_io_in_psum = PE_Array_7_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_15_clock = clock;
  assign PE_Array_8_15_reset = reset;
  assign PE_Array_8_15_io_in_activate = PE_Array_8_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_15_io_in_weight = PE_Array_7_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_15_io_in_psum = PE_Array_7_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_0_clock = clock;
  assign PE_Array_9_0_reset = reset;
  assign PE_Array_9_0_io_in_activate = io_activate_9; // @[DataPath.scala 11:26]
  assign PE_Array_9_0_io_in_weight = PE_Array_8_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_0_io_in_psum = PE_Array_8_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_1_clock = clock;
  assign PE_Array_9_1_reset = reset;
  assign PE_Array_9_1_io_in_activate = PE_Array_9_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_1_io_in_weight = PE_Array_8_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_1_io_in_psum = PE_Array_8_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_2_clock = clock;
  assign PE_Array_9_2_reset = reset;
  assign PE_Array_9_2_io_in_activate = PE_Array_9_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_2_io_in_weight = PE_Array_8_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_2_io_in_psum = PE_Array_8_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_3_clock = clock;
  assign PE_Array_9_3_reset = reset;
  assign PE_Array_9_3_io_in_activate = PE_Array_9_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_3_io_in_weight = PE_Array_8_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_3_io_in_psum = PE_Array_8_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_4_clock = clock;
  assign PE_Array_9_4_reset = reset;
  assign PE_Array_9_4_io_in_activate = PE_Array_9_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_4_io_in_weight = PE_Array_8_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_4_io_in_psum = PE_Array_8_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_5_clock = clock;
  assign PE_Array_9_5_reset = reset;
  assign PE_Array_9_5_io_in_activate = PE_Array_9_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_5_io_in_weight = PE_Array_8_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_5_io_in_psum = PE_Array_8_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_6_clock = clock;
  assign PE_Array_9_6_reset = reset;
  assign PE_Array_9_6_io_in_activate = PE_Array_9_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_6_io_in_weight = PE_Array_8_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_6_io_in_psum = PE_Array_8_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_7_clock = clock;
  assign PE_Array_9_7_reset = reset;
  assign PE_Array_9_7_io_in_activate = PE_Array_9_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_7_io_in_weight = PE_Array_8_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_7_io_in_psum = PE_Array_8_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_8_clock = clock;
  assign PE_Array_9_8_reset = reset;
  assign PE_Array_9_8_io_in_activate = PE_Array_9_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_8_io_in_weight = PE_Array_8_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_8_io_in_psum = PE_Array_8_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_9_clock = clock;
  assign PE_Array_9_9_reset = reset;
  assign PE_Array_9_9_io_in_activate = PE_Array_9_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_9_io_in_weight = PE_Array_8_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_9_io_in_psum = PE_Array_8_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_10_clock = clock;
  assign PE_Array_9_10_reset = reset;
  assign PE_Array_9_10_io_in_activate = PE_Array_9_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_10_io_in_weight = PE_Array_8_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_10_io_in_psum = PE_Array_8_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_11_clock = clock;
  assign PE_Array_9_11_reset = reset;
  assign PE_Array_9_11_io_in_activate = PE_Array_9_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_11_io_in_weight = PE_Array_8_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_11_io_in_psum = PE_Array_8_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_12_clock = clock;
  assign PE_Array_9_12_reset = reset;
  assign PE_Array_9_12_io_in_activate = PE_Array_9_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_12_io_in_weight = PE_Array_8_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_12_io_in_psum = PE_Array_8_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_13_clock = clock;
  assign PE_Array_9_13_reset = reset;
  assign PE_Array_9_13_io_in_activate = PE_Array_9_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_13_io_in_weight = PE_Array_8_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_13_io_in_psum = PE_Array_8_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_14_clock = clock;
  assign PE_Array_9_14_reset = reset;
  assign PE_Array_9_14_io_in_activate = PE_Array_9_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_14_io_in_weight = PE_Array_8_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_14_io_in_psum = PE_Array_8_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_15_clock = clock;
  assign PE_Array_9_15_reset = reset;
  assign PE_Array_9_15_io_in_activate = PE_Array_9_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_15_io_in_weight = PE_Array_8_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_15_io_in_psum = PE_Array_8_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_0_clock = clock;
  assign PE_Array_10_0_reset = reset;
  assign PE_Array_10_0_io_in_activate = io_activate_10; // @[DataPath.scala 11:26]
  assign PE_Array_10_0_io_in_weight = PE_Array_9_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_0_io_in_psum = PE_Array_9_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_1_clock = clock;
  assign PE_Array_10_1_reset = reset;
  assign PE_Array_10_1_io_in_activate = PE_Array_10_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_1_io_in_weight = PE_Array_9_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_1_io_in_psum = PE_Array_9_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_2_clock = clock;
  assign PE_Array_10_2_reset = reset;
  assign PE_Array_10_2_io_in_activate = PE_Array_10_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_2_io_in_weight = PE_Array_9_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_2_io_in_psum = PE_Array_9_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_3_clock = clock;
  assign PE_Array_10_3_reset = reset;
  assign PE_Array_10_3_io_in_activate = PE_Array_10_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_3_io_in_weight = PE_Array_9_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_3_io_in_psum = PE_Array_9_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_4_clock = clock;
  assign PE_Array_10_4_reset = reset;
  assign PE_Array_10_4_io_in_activate = PE_Array_10_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_4_io_in_weight = PE_Array_9_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_4_io_in_psum = PE_Array_9_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_5_clock = clock;
  assign PE_Array_10_5_reset = reset;
  assign PE_Array_10_5_io_in_activate = PE_Array_10_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_5_io_in_weight = PE_Array_9_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_5_io_in_psum = PE_Array_9_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_6_clock = clock;
  assign PE_Array_10_6_reset = reset;
  assign PE_Array_10_6_io_in_activate = PE_Array_10_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_6_io_in_weight = PE_Array_9_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_6_io_in_psum = PE_Array_9_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_7_clock = clock;
  assign PE_Array_10_7_reset = reset;
  assign PE_Array_10_7_io_in_activate = PE_Array_10_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_7_io_in_weight = PE_Array_9_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_7_io_in_psum = PE_Array_9_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_8_clock = clock;
  assign PE_Array_10_8_reset = reset;
  assign PE_Array_10_8_io_in_activate = PE_Array_10_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_8_io_in_weight = PE_Array_9_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_8_io_in_psum = PE_Array_9_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_9_clock = clock;
  assign PE_Array_10_9_reset = reset;
  assign PE_Array_10_9_io_in_activate = PE_Array_10_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_9_io_in_weight = PE_Array_9_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_9_io_in_psum = PE_Array_9_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_10_clock = clock;
  assign PE_Array_10_10_reset = reset;
  assign PE_Array_10_10_io_in_activate = PE_Array_10_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_10_io_in_weight = PE_Array_9_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_10_io_in_psum = PE_Array_9_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_11_clock = clock;
  assign PE_Array_10_11_reset = reset;
  assign PE_Array_10_11_io_in_activate = PE_Array_10_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_11_io_in_weight = PE_Array_9_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_11_io_in_psum = PE_Array_9_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_12_clock = clock;
  assign PE_Array_10_12_reset = reset;
  assign PE_Array_10_12_io_in_activate = PE_Array_10_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_12_io_in_weight = PE_Array_9_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_12_io_in_psum = PE_Array_9_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_13_clock = clock;
  assign PE_Array_10_13_reset = reset;
  assign PE_Array_10_13_io_in_activate = PE_Array_10_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_13_io_in_weight = PE_Array_9_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_13_io_in_psum = PE_Array_9_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_14_clock = clock;
  assign PE_Array_10_14_reset = reset;
  assign PE_Array_10_14_io_in_activate = PE_Array_10_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_14_io_in_weight = PE_Array_9_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_14_io_in_psum = PE_Array_9_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_15_clock = clock;
  assign PE_Array_10_15_reset = reset;
  assign PE_Array_10_15_io_in_activate = PE_Array_10_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_15_io_in_weight = PE_Array_9_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_15_io_in_psum = PE_Array_9_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_0_clock = clock;
  assign PE_Array_11_0_reset = reset;
  assign PE_Array_11_0_io_in_activate = io_activate_11; // @[DataPath.scala 11:26]
  assign PE_Array_11_0_io_in_weight = PE_Array_10_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_0_io_in_psum = PE_Array_10_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_1_clock = clock;
  assign PE_Array_11_1_reset = reset;
  assign PE_Array_11_1_io_in_activate = PE_Array_11_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_1_io_in_weight = PE_Array_10_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_1_io_in_psum = PE_Array_10_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_2_clock = clock;
  assign PE_Array_11_2_reset = reset;
  assign PE_Array_11_2_io_in_activate = PE_Array_11_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_2_io_in_weight = PE_Array_10_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_2_io_in_psum = PE_Array_10_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_3_clock = clock;
  assign PE_Array_11_3_reset = reset;
  assign PE_Array_11_3_io_in_activate = PE_Array_11_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_3_io_in_weight = PE_Array_10_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_3_io_in_psum = PE_Array_10_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_4_clock = clock;
  assign PE_Array_11_4_reset = reset;
  assign PE_Array_11_4_io_in_activate = PE_Array_11_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_4_io_in_weight = PE_Array_10_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_4_io_in_psum = PE_Array_10_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_5_clock = clock;
  assign PE_Array_11_5_reset = reset;
  assign PE_Array_11_5_io_in_activate = PE_Array_11_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_5_io_in_weight = PE_Array_10_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_5_io_in_psum = PE_Array_10_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_6_clock = clock;
  assign PE_Array_11_6_reset = reset;
  assign PE_Array_11_6_io_in_activate = PE_Array_11_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_6_io_in_weight = PE_Array_10_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_6_io_in_psum = PE_Array_10_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_7_clock = clock;
  assign PE_Array_11_7_reset = reset;
  assign PE_Array_11_7_io_in_activate = PE_Array_11_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_7_io_in_weight = PE_Array_10_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_7_io_in_psum = PE_Array_10_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_8_clock = clock;
  assign PE_Array_11_8_reset = reset;
  assign PE_Array_11_8_io_in_activate = PE_Array_11_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_8_io_in_weight = PE_Array_10_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_8_io_in_psum = PE_Array_10_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_9_clock = clock;
  assign PE_Array_11_9_reset = reset;
  assign PE_Array_11_9_io_in_activate = PE_Array_11_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_9_io_in_weight = PE_Array_10_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_9_io_in_psum = PE_Array_10_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_10_clock = clock;
  assign PE_Array_11_10_reset = reset;
  assign PE_Array_11_10_io_in_activate = PE_Array_11_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_10_io_in_weight = PE_Array_10_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_10_io_in_psum = PE_Array_10_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_11_clock = clock;
  assign PE_Array_11_11_reset = reset;
  assign PE_Array_11_11_io_in_activate = PE_Array_11_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_11_io_in_weight = PE_Array_10_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_11_io_in_psum = PE_Array_10_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_12_clock = clock;
  assign PE_Array_11_12_reset = reset;
  assign PE_Array_11_12_io_in_activate = PE_Array_11_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_12_io_in_weight = PE_Array_10_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_12_io_in_psum = PE_Array_10_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_13_clock = clock;
  assign PE_Array_11_13_reset = reset;
  assign PE_Array_11_13_io_in_activate = PE_Array_11_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_13_io_in_weight = PE_Array_10_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_13_io_in_psum = PE_Array_10_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_14_clock = clock;
  assign PE_Array_11_14_reset = reset;
  assign PE_Array_11_14_io_in_activate = PE_Array_11_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_14_io_in_weight = PE_Array_10_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_14_io_in_psum = PE_Array_10_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_15_clock = clock;
  assign PE_Array_11_15_reset = reset;
  assign PE_Array_11_15_io_in_activate = PE_Array_11_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_15_io_in_weight = PE_Array_10_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_15_io_in_psum = PE_Array_10_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_0_clock = clock;
  assign PE_Array_12_0_reset = reset;
  assign PE_Array_12_0_io_in_activate = io_activate_12; // @[DataPath.scala 11:26]
  assign PE_Array_12_0_io_in_weight = PE_Array_11_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_0_io_in_psum = PE_Array_11_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_1_clock = clock;
  assign PE_Array_12_1_reset = reset;
  assign PE_Array_12_1_io_in_activate = PE_Array_12_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_1_io_in_weight = PE_Array_11_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_1_io_in_psum = PE_Array_11_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_2_clock = clock;
  assign PE_Array_12_2_reset = reset;
  assign PE_Array_12_2_io_in_activate = PE_Array_12_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_2_io_in_weight = PE_Array_11_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_2_io_in_psum = PE_Array_11_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_3_clock = clock;
  assign PE_Array_12_3_reset = reset;
  assign PE_Array_12_3_io_in_activate = PE_Array_12_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_3_io_in_weight = PE_Array_11_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_3_io_in_psum = PE_Array_11_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_4_clock = clock;
  assign PE_Array_12_4_reset = reset;
  assign PE_Array_12_4_io_in_activate = PE_Array_12_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_4_io_in_weight = PE_Array_11_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_4_io_in_psum = PE_Array_11_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_5_clock = clock;
  assign PE_Array_12_5_reset = reset;
  assign PE_Array_12_5_io_in_activate = PE_Array_12_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_5_io_in_weight = PE_Array_11_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_5_io_in_psum = PE_Array_11_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_6_clock = clock;
  assign PE_Array_12_6_reset = reset;
  assign PE_Array_12_6_io_in_activate = PE_Array_12_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_6_io_in_weight = PE_Array_11_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_6_io_in_psum = PE_Array_11_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_7_clock = clock;
  assign PE_Array_12_7_reset = reset;
  assign PE_Array_12_7_io_in_activate = PE_Array_12_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_7_io_in_weight = PE_Array_11_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_7_io_in_psum = PE_Array_11_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_8_clock = clock;
  assign PE_Array_12_8_reset = reset;
  assign PE_Array_12_8_io_in_activate = PE_Array_12_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_8_io_in_weight = PE_Array_11_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_8_io_in_psum = PE_Array_11_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_9_clock = clock;
  assign PE_Array_12_9_reset = reset;
  assign PE_Array_12_9_io_in_activate = PE_Array_12_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_9_io_in_weight = PE_Array_11_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_9_io_in_psum = PE_Array_11_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_10_clock = clock;
  assign PE_Array_12_10_reset = reset;
  assign PE_Array_12_10_io_in_activate = PE_Array_12_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_10_io_in_weight = PE_Array_11_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_10_io_in_psum = PE_Array_11_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_11_clock = clock;
  assign PE_Array_12_11_reset = reset;
  assign PE_Array_12_11_io_in_activate = PE_Array_12_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_11_io_in_weight = PE_Array_11_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_11_io_in_psum = PE_Array_11_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_12_clock = clock;
  assign PE_Array_12_12_reset = reset;
  assign PE_Array_12_12_io_in_activate = PE_Array_12_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_12_io_in_weight = PE_Array_11_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_12_io_in_psum = PE_Array_11_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_13_clock = clock;
  assign PE_Array_12_13_reset = reset;
  assign PE_Array_12_13_io_in_activate = PE_Array_12_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_13_io_in_weight = PE_Array_11_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_13_io_in_psum = PE_Array_11_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_14_clock = clock;
  assign PE_Array_12_14_reset = reset;
  assign PE_Array_12_14_io_in_activate = PE_Array_12_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_14_io_in_weight = PE_Array_11_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_14_io_in_psum = PE_Array_11_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_15_clock = clock;
  assign PE_Array_12_15_reset = reset;
  assign PE_Array_12_15_io_in_activate = PE_Array_12_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_15_io_in_weight = PE_Array_11_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_15_io_in_psum = PE_Array_11_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_0_clock = clock;
  assign PE_Array_13_0_reset = reset;
  assign PE_Array_13_0_io_in_activate = io_activate_13; // @[DataPath.scala 11:26]
  assign PE_Array_13_0_io_in_weight = PE_Array_12_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_0_io_in_psum = PE_Array_12_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_1_clock = clock;
  assign PE_Array_13_1_reset = reset;
  assign PE_Array_13_1_io_in_activate = PE_Array_13_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_1_io_in_weight = PE_Array_12_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_1_io_in_psum = PE_Array_12_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_2_clock = clock;
  assign PE_Array_13_2_reset = reset;
  assign PE_Array_13_2_io_in_activate = PE_Array_13_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_2_io_in_weight = PE_Array_12_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_2_io_in_psum = PE_Array_12_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_3_clock = clock;
  assign PE_Array_13_3_reset = reset;
  assign PE_Array_13_3_io_in_activate = PE_Array_13_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_3_io_in_weight = PE_Array_12_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_3_io_in_psum = PE_Array_12_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_4_clock = clock;
  assign PE_Array_13_4_reset = reset;
  assign PE_Array_13_4_io_in_activate = PE_Array_13_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_4_io_in_weight = PE_Array_12_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_4_io_in_psum = PE_Array_12_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_5_clock = clock;
  assign PE_Array_13_5_reset = reset;
  assign PE_Array_13_5_io_in_activate = PE_Array_13_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_5_io_in_weight = PE_Array_12_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_5_io_in_psum = PE_Array_12_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_6_clock = clock;
  assign PE_Array_13_6_reset = reset;
  assign PE_Array_13_6_io_in_activate = PE_Array_13_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_6_io_in_weight = PE_Array_12_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_6_io_in_psum = PE_Array_12_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_7_clock = clock;
  assign PE_Array_13_7_reset = reset;
  assign PE_Array_13_7_io_in_activate = PE_Array_13_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_7_io_in_weight = PE_Array_12_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_7_io_in_psum = PE_Array_12_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_8_clock = clock;
  assign PE_Array_13_8_reset = reset;
  assign PE_Array_13_8_io_in_activate = PE_Array_13_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_8_io_in_weight = PE_Array_12_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_8_io_in_psum = PE_Array_12_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_9_clock = clock;
  assign PE_Array_13_9_reset = reset;
  assign PE_Array_13_9_io_in_activate = PE_Array_13_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_9_io_in_weight = PE_Array_12_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_9_io_in_psum = PE_Array_12_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_10_clock = clock;
  assign PE_Array_13_10_reset = reset;
  assign PE_Array_13_10_io_in_activate = PE_Array_13_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_10_io_in_weight = PE_Array_12_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_10_io_in_psum = PE_Array_12_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_11_clock = clock;
  assign PE_Array_13_11_reset = reset;
  assign PE_Array_13_11_io_in_activate = PE_Array_13_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_11_io_in_weight = PE_Array_12_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_11_io_in_psum = PE_Array_12_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_12_clock = clock;
  assign PE_Array_13_12_reset = reset;
  assign PE_Array_13_12_io_in_activate = PE_Array_13_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_12_io_in_weight = PE_Array_12_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_12_io_in_psum = PE_Array_12_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_13_clock = clock;
  assign PE_Array_13_13_reset = reset;
  assign PE_Array_13_13_io_in_activate = PE_Array_13_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_13_io_in_weight = PE_Array_12_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_13_io_in_psum = PE_Array_12_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_14_clock = clock;
  assign PE_Array_13_14_reset = reset;
  assign PE_Array_13_14_io_in_activate = PE_Array_13_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_14_io_in_weight = PE_Array_12_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_14_io_in_psum = PE_Array_12_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_15_clock = clock;
  assign PE_Array_13_15_reset = reset;
  assign PE_Array_13_15_io_in_activate = PE_Array_13_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_15_io_in_weight = PE_Array_12_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_15_io_in_psum = PE_Array_12_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_0_clock = clock;
  assign PE_Array_14_0_reset = reset;
  assign PE_Array_14_0_io_in_activate = io_activate_14; // @[DataPath.scala 11:26]
  assign PE_Array_14_0_io_in_weight = PE_Array_13_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_0_io_in_psum = PE_Array_13_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_1_clock = clock;
  assign PE_Array_14_1_reset = reset;
  assign PE_Array_14_1_io_in_activate = PE_Array_14_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_1_io_in_weight = PE_Array_13_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_1_io_in_psum = PE_Array_13_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_2_clock = clock;
  assign PE_Array_14_2_reset = reset;
  assign PE_Array_14_2_io_in_activate = PE_Array_14_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_2_io_in_weight = PE_Array_13_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_2_io_in_psum = PE_Array_13_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_3_clock = clock;
  assign PE_Array_14_3_reset = reset;
  assign PE_Array_14_3_io_in_activate = PE_Array_14_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_3_io_in_weight = PE_Array_13_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_3_io_in_psum = PE_Array_13_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_4_clock = clock;
  assign PE_Array_14_4_reset = reset;
  assign PE_Array_14_4_io_in_activate = PE_Array_14_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_4_io_in_weight = PE_Array_13_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_4_io_in_psum = PE_Array_13_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_5_clock = clock;
  assign PE_Array_14_5_reset = reset;
  assign PE_Array_14_5_io_in_activate = PE_Array_14_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_5_io_in_weight = PE_Array_13_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_5_io_in_psum = PE_Array_13_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_6_clock = clock;
  assign PE_Array_14_6_reset = reset;
  assign PE_Array_14_6_io_in_activate = PE_Array_14_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_6_io_in_weight = PE_Array_13_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_6_io_in_psum = PE_Array_13_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_7_clock = clock;
  assign PE_Array_14_7_reset = reset;
  assign PE_Array_14_7_io_in_activate = PE_Array_14_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_7_io_in_weight = PE_Array_13_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_7_io_in_psum = PE_Array_13_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_8_clock = clock;
  assign PE_Array_14_8_reset = reset;
  assign PE_Array_14_8_io_in_activate = PE_Array_14_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_8_io_in_weight = PE_Array_13_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_8_io_in_psum = PE_Array_13_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_9_clock = clock;
  assign PE_Array_14_9_reset = reset;
  assign PE_Array_14_9_io_in_activate = PE_Array_14_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_9_io_in_weight = PE_Array_13_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_9_io_in_psum = PE_Array_13_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_10_clock = clock;
  assign PE_Array_14_10_reset = reset;
  assign PE_Array_14_10_io_in_activate = PE_Array_14_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_10_io_in_weight = PE_Array_13_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_10_io_in_psum = PE_Array_13_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_11_clock = clock;
  assign PE_Array_14_11_reset = reset;
  assign PE_Array_14_11_io_in_activate = PE_Array_14_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_11_io_in_weight = PE_Array_13_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_11_io_in_psum = PE_Array_13_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_12_clock = clock;
  assign PE_Array_14_12_reset = reset;
  assign PE_Array_14_12_io_in_activate = PE_Array_14_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_12_io_in_weight = PE_Array_13_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_12_io_in_psum = PE_Array_13_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_13_clock = clock;
  assign PE_Array_14_13_reset = reset;
  assign PE_Array_14_13_io_in_activate = PE_Array_14_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_13_io_in_weight = PE_Array_13_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_13_io_in_psum = PE_Array_13_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_14_clock = clock;
  assign PE_Array_14_14_reset = reset;
  assign PE_Array_14_14_io_in_activate = PE_Array_14_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_14_io_in_weight = PE_Array_13_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_14_io_in_psum = PE_Array_13_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_15_clock = clock;
  assign PE_Array_14_15_reset = reset;
  assign PE_Array_14_15_io_in_activate = PE_Array_14_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_15_io_in_weight = PE_Array_13_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_15_io_in_psum = PE_Array_13_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_0_clock = clock;
  assign PE_Array_15_0_reset = reset;
  assign PE_Array_15_0_io_in_activate = io_activate_15; // @[DataPath.scala 11:26]
  assign PE_Array_15_0_io_in_weight = PE_Array_14_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_0_io_in_psum = PE_Array_14_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_1_clock = clock;
  assign PE_Array_15_1_reset = reset;
  assign PE_Array_15_1_io_in_activate = PE_Array_15_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_1_io_in_weight = PE_Array_14_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_1_io_in_psum = PE_Array_14_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_2_clock = clock;
  assign PE_Array_15_2_reset = reset;
  assign PE_Array_15_2_io_in_activate = PE_Array_15_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_2_io_in_weight = PE_Array_14_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_2_io_in_psum = PE_Array_14_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_3_clock = clock;
  assign PE_Array_15_3_reset = reset;
  assign PE_Array_15_3_io_in_activate = PE_Array_15_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_3_io_in_weight = PE_Array_14_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_3_io_in_psum = PE_Array_14_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_4_clock = clock;
  assign PE_Array_15_4_reset = reset;
  assign PE_Array_15_4_io_in_activate = PE_Array_15_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_4_io_in_weight = PE_Array_14_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_4_io_in_psum = PE_Array_14_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_5_clock = clock;
  assign PE_Array_15_5_reset = reset;
  assign PE_Array_15_5_io_in_activate = PE_Array_15_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_5_io_in_weight = PE_Array_14_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_5_io_in_psum = PE_Array_14_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_6_clock = clock;
  assign PE_Array_15_6_reset = reset;
  assign PE_Array_15_6_io_in_activate = PE_Array_15_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_6_io_in_weight = PE_Array_14_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_6_io_in_psum = PE_Array_14_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_7_clock = clock;
  assign PE_Array_15_7_reset = reset;
  assign PE_Array_15_7_io_in_activate = PE_Array_15_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_7_io_in_weight = PE_Array_14_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_7_io_in_psum = PE_Array_14_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_8_clock = clock;
  assign PE_Array_15_8_reset = reset;
  assign PE_Array_15_8_io_in_activate = PE_Array_15_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_8_io_in_weight = PE_Array_14_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_8_io_in_psum = PE_Array_14_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_9_clock = clock;
  assign PE_Array_15_9_reset = reset;
  assign PE_Array_15_9_io_in_activate = PE_Array_15_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_9_io_in_weight = PE_Array_14_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_9_io_in_psum = PE_Array_14_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_10_clock = clock;
  assign PE_Array_15_10_reset = reset;
  assign PE_Array_15_10_io_in_activate = PE_Array_15_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_10_io_in_weight = PE_Array_14_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_10_io_in_psum = PE_Array_14_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_11_clock = clock;
  assign PE_Array_15_11_reset = reset;
  assign PE_Array_15_11_io_in_activate = PE_Array_15_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_11_io_in_weight = PE_Array_14_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_11_io_in_psum = PE_Array_14_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_12_clock = clock;
  assign PE_Array_15_12_reset = reset;
  assign PE_Array_15_12_io_in_activate = PE_Array_15_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_12_io_in_weight = PE_Array_14_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_12_io_in_psum = PE_Array_14_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_13_clock = clock;
  assign PE_Array_15_13_reset = reset;
  assign PE_Array_15_13_io_in_activate = PE_Array_15_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_13_io_in_weight = PE_Array_14_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_13_io_in_psum = PE_Array_14_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_14_clock = clock;
  assign PE_Array_15_14_reset = reset;
  assign PE_Array_15_14_io_in_activate = PE_Array_15_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_14_io_in_weight = PE_Array_14_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_14_io_in_psum = PE_Array_14_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_15_clock = clock;
  assign PE_Array_15_15_reset = reset;
  assign PE_Array_15_15_io_in_activate = PE_Array_15_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_15_io_in_weight = PE_Array_14_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_15_io_in_psum = PE_Array_14_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  always @(posedge clock) begin
    if (reset) begin // @[Systolic_Array.scala 52:29]
      flow_counter <= 6'h0; // @[Systolic_Array.scala 52:29]
    end else if (io_flow & flow_counter < 6'h2e) begin // @[Systolic_Array.scala 56:58]
      flow_counter <= _flow_counter_T_1; // @[Systolic_Array.scala 57:18]
    end else if (flow_counter == 6'h2e) begin // @[Systolic_Array.scala 58:53]
      flow_counter <= 6'h0; // @[Systolic_Array.scala 59:18]
    end
    if (reset) begin // @[Systolic_Array.scala 53:26]
      valid_reg <= 16'h0; // @[Systolic_Array.scala 53:26]
    end else if (io_flow & 6'hf <= flow_counter & flow_counter < 6'h1f) begin // @[Systolic_Array.scala 65:96]
      valid_reg <= _valid_reg_T_1; // @[Systolic_Array.scala 66:15]
    end else if (io_flow & flow_counter >= 6'h1f) begin // @[Systolic_Array.scala 67:65]
      valid_reg <= _valid_reg_T_3; // @[Systolic_Array.scala 68:15]
    end else begin
      valid_reg <= 16'h0; // @[Systolic_Array.scala 70:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flow_counter = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
