module basic_PE(
  input         clock,
  input         reset,
  input  [7:0]  io_in_activate,
  input  [7:0]  io_in_weight,
  input  [15:0] io_in_psum,
  input         io_in_flow,
  input         io_in_shift,
  output [7:0]  io_out_activate,
  output [7:0]  io_out_weight,
  output [15:0] io_out_psum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] Activation_Reg; // @[basic_PE.scala 17:31]
  reg [7:0] Weight_Reg; // @[basic_PE.scala 18:27]
  reg [15:0] PSum_Reg; // @[basic_PE.scala 19:25]
  wire [15:0] _io_out_psum_T = Activation_Reg * Weight_Reg; // @[basic_PE.scala 47:33]
  assign io_out_activate = Activation_Reg; // @[basic_PE.scala 45:19]
  assign io_out_weight = Weight_Reg; // @[basic_PE.scala 46:17]
  assign io_out_psum = _io_out_psum_T + PSum_Reg; // @[basic_PE.scala 47:46]
  always @(posedge clock) begin
    if (reset) begin // @[basic_PE.scala 17:31]
      Activation_Reg <= 8'h0; // @[basic_PE.scala 17:31]
    end else if (io_in_flow) begin // @[basic_PE.scala 22:20]
      Activation_Reg <= io_in_activate; // @[basic_PE.scala 23:20]
    end
    if (reset) begin // @[basic_PE.scala 18:27]
      Weight_Reg <= 8'h0; // @[basic_PE.scala 18:27]
    end else if (io_in_shift) begin // @[basic_PE.scala 38:21]
      Weight_Reg <= io_in_weight; // @[basic_PE.scala 39:16]
    end
    if (reset) begin // @[basic_PE.scala 19:25]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 19:25]
    end else if (io_in_shift) begin // @[basic_PE.scala 29:21]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 30:14]
    end else if (io_in_flow) begin // @[basic_PE.scala 31:26]
      PSum_Reg <= io_in_psum; // @[basic_PE.scala 32:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Activation_Reg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  Weight_Reg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  PSum_Reg = _RAND_2[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Systolic_Array(
  input         clock,
  input         reset,
  input  [7:0]  io_activate_0,
  input  [7:0]  io_activate_1,
  input  [7:0]  io_activate_2,
  input  [7:0]  io_activate_3,
  input  [7:0]  io_activate_4,
  input  [7:0]  io_activate_5,
  input  [7:0]  io_activate_6,
  input  [7:0]  io_activate_7,
  input  [7:0]  io_activate_8,
  input  [7:0]  io_activate_9,
  input  [7:0]  io_activate_10,
  input  [7:0]  io_activate_11,
  input  [7:0]  io_activate_12,
  input  [7:0]  io_activate_13,
  input  [7:0]  io_activate_14,
  input  [7:0]  io_activate_15,
  input  [7:0]  io_activate_16,
  input  [7:0]  io_activate_17,
  input  [7:0]  io_activate_18,
  input  [7:0]  io_activate_19,
  input  [7:0]  io_activate_20,
  input  [7:0]  io_activate_21,
  input  [7:0]  io_activate_22,
  input  [7:0]  io_activate_23,
  input  [7:0]  io_activate_24,
  input  [7:0]  io_activate_25,
  input  [7:0]  io_activate_26,
  input  [7:0]  io_activate_27,
  input  [7:0]  io_activate_28,
  input  [7:0]  io_activate_29,
  input  [7:0]  io_activate_30,
  input  [7:0]  io_activate_31,
  input  [7:0]  io_weight_0,
  input  [7:0]  io_weight_1,
  input  [7:0]  io_weight_2,
  input  [7:0]  io_weight_3,
  input  [7:0]  io_weight_4,
  input  [7:0]  io_weight_5,
  input  [7:0]  io_weight_6,
  input  [7:0]  io_weight_7,
  input  [7:0]  io_weight_8,
  input  [7:0]  io_weight_9,
  input  [7:0]  io_weight_10,
  input  [7:0]  io_weight_11,
  input  [7:0]  io_weight_12,
  input  [7:0]  io_weight_13,
  input  [7:0]  io_weight_14,
  input  [7:0]  io_weight_15,
  input  [7:0]  io_weight_16,
  input  [7:0]  io_weight_17,
  input  [7:0]  io_weight_18,
  input  [7:0]  io_weight_19,
  input  [7:0]  io_weight_20,
  input  [7:0]  io_weight_21,
  input  [7:0]  io_weight_22,
  input  [7:0]  io_weight_23,
  input  [7:0]  io_weight_24,
  input  [7:0]  io_weight_25,
  input  [7:0]  io_weight_26,
  input  [7:0]  io_weight_27,
  input  [7:0]  io_weight_28,
  input  [7:0]  io_weight_29,
  input  [7:0]  io_weight_30,
  input  [7:0]  io_weight_31,
  input         io_flow,
  input         io_shift,
  output [15:0] io_psum_0,
  output [15:0] io_psum_1,
  output [15:0] io_psum_2,
  output [15:0] io_psum_3,
  output [15:0] io_psum_4,
  output [15:0] io_psum_5,
  output [15:0] io_psum_6,
  output [15:0] io_psum_7,
  output [15:0] io_psum_8,
  output [15:0] io_psum_9,
  output [15:0] io_psum_10,
  output [15:0] io_psum_11,
  output [15:0] io_psum_12,
  output [15:0] io_psum_13,
  output [15:0] io_psum_14,
  output [15:0] io_psum_15,
  output [15:0] io_psum_16,
  output [15:0] io_psum_17,
  output [15:0] io_psum_18,
  output [15:0] io_psum_19,
  output [15:0] io_psum_20,
  output [15:0] io_psum_21,
  output [15:0] io_psum_22,
  output [15:0] io_psum_23,
  output [15:0] io_psum_24,
  output [15:0] io_psum_25,
  output [15:0] io_psum_26,
  output [15:0] io_psum_27,
  output [15:0] io_psum_28,
  output [15:0] io_psum_29,
  output [15:0] io_psum_30,
  output [15:0] io_psum_31,
  output        io_valid_0,
  output        io_valid_1,
  output        io_valid_2,
  output        io_valid_3,
  output        io_valid_4,
  output        io_valid_5,
  output        io_valid_6,
  output        io_valid_7,
  output        io_valid_8,
  output        io_valid_9,
  output        io_valid_10,
  output        io_valid_11,
  output        io_valid_12,
  output        io_valid_13,
  output        io_valid_14,
  output        io_valid_15,
  output        io_valid_16,
  output        io_valid_17,
  output        io_valid_18,
  output        io_valid_19,
  output        io_valid_20,
  output        io_valid_21,
  output        io_valid_22,
  output        io_valid_23,
  output        io_valid_24,
  output        io_valid_25,
  output        io_valid_26,
  output        io_valid_27,
  output        io_valid_28,
  output        io_valid_29,
  output        io_valid_30,
  output        io_valid_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  PE_Array_0_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_8_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_8_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_8_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_9_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_9_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_9_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_10_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_10_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_10_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_11_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_11_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_11_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_12_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_12_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_12_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_13_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_13_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_13_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_14_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_14_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_14_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_15_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_15_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_15_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_16_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_16_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_16_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_17_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_17_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_17_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_18_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_18_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_18_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_19_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_19_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_19_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_20_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_20_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_20_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_21_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_21_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_21_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_22_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_22_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_22_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_23_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_23_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_23_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_24_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_24_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_24_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_25_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_25_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_25_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_26_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_26_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_26_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_27_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_27_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_27_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_28_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_28_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_28_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_29_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_29_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_29_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_30_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_30_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_30_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_8_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_8_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_8_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_8_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_8_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_8_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_8_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_8_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_8_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_8_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_9_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_9_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_9_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_9_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_9_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_9_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_9_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_9_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_9_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_9_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_10_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_10_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_10_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_10_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_10_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_10_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_10_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_10_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_10_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_10_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_11_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_11_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_11_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_11_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_11_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_11_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_11_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_11_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_11_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_11_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_12_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_12_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_12_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_12_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_12_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_12_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_12_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_12_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_12_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_12_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_13_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_13_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_13_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_13_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_13_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_13_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_13_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_13_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_13_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_13_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_14_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_14_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_14_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_14_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_14_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_14_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_14_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_14_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_14_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_14_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_15_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_15_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_15_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_15_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_15_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_15_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_15_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_15_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_15_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_15_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_16_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_16_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_16_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_16_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_16_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_16_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_16_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_16_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_16_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_16_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_17_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_17_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_17_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_17_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_17_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_17_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_17_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_17_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_17_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_17_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_18_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_18_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_18_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_18_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_18_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_18_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_18_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_18_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_18_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_18_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_19_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_19_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_19_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_19_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_19_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_19_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_19_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_19_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_19_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_19_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_20_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_20_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_20_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_20_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_20_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_20_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_20_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_20_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_20_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_20_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_21_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_21_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_21_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_21_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_21_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_21_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_21_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_21_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_21_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_21_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_22_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_22_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_22_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_22_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_22_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_22_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_22_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_22_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_22_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_22_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_23_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_23_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_23_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_23_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_23_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_23_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_23_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_23_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_23_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_23_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_24_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_24_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_24_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_24_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_24_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_24_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_24_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_24_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_24_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_24_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_25_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_25_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_25_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_25_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_25_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_25_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_25_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_25_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_25_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_25_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_26_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_26_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_26_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_26_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_26_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_26_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_26_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_26_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_26_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_26_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_27_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_27_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_27_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_27_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_27_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_27_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_27_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_27_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_27_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_27_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_28_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_28_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_28_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_28_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_28_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_28_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_28_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_28_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_28_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_28_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_29_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_29_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_29_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_29_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_29_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_29_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_29_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_29_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_29_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_29_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_30_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_30_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_30_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_30_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_30_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_30_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_30_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_30_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_30_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_30_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_31_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_31_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_31_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_31_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_31_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_31_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_31_31_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_31_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_31_31_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_31_31_io_out_psum; // @[Systolic_Array.scala 19:62]
  reg [6:0] flow_counter; // @[Systolic_Array.scala 52:29]
  reg [31:0] valid_reg; // @[Systolic_Array.scala 53:26]
  wire [6:0] _flow_counter_T_1 = flow_counter + 7'h1; // @[Systolic_Array.scala 57:34]
  wire [31:0] _valid_reg_T_1 = {valid_reg[30:0],1'h1}; // @[Cat.scala 33:92]
  wire [31:0] _valid_reg_T_3 = {valid_reg[30:0],1'h0}; // @[Cat.scala 33:92]
  basic_PE PE_Array_0_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_0_clock),
    .reset(PE_Array_0_0_reset),
    .io_in_activate(PE_Array_0_0_io_in_activate),
    .io_in_weight(PE_Array_0_0_io_in_weight),
    .io_in_psum(PE_Array_0_0_io_in_psum),
    .io_in_flow(PE_Array_0_0_io_in_flow),
    .io_in_shift(PE_Array_0_0_io_in_shift),
    .io_out_activate(PE_Array_0_0_io_out_activate),
    .io_out_weight(PE_Array_0_0_io_out_weight),
    .io_out_psum(PE_Array_0_0_io_out_psum)
  );
  basic_PE PE_Array_0_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_1_clock),
    .reset(PE_Array_0_1_reset),
    .io_in_activate(PE_Array_0_1_io_in_activate),
    .io_in_weight(PE_Array_0_1_io_in_weight),
    .io_in_psum(PE_Array_0_1_io_in_psum),
    .io_in_flow(PE_Array_0_1_io_in_flow),
    .io_in_shift(PE_Array_0_1_io_in_shift),
    .io_out_activate(PE_Array_0_1_io_out_activate),
    .io_out_weight(PE_Array_0_1_io_out_weight),
    .io_out_psum(PE_Array_0_1_io_out_psum)
  );
  basic_PE PE_Array_0_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_2_clock),
    .reset(PE_Array_0_2_reset),
    .io_in_activate(PE_Array_0_2_io_in_activate),
    .io_in_weight(PE_Array_0_2_io_in_weight),
    .io_in_psum(PE_Array_0_2_io_in_psum),
    .io_in_flow(PE_Array_0_2_io_in_flow),
    .io_in_shift(PE_Array_0_2_io_in_shift),
    .io_out_activate(PE_Array_0_2_io_out_activate),
    .io_out_weight(PE_Array_0_2_io_out_weight),
    .io_out_psum(PE_Array_0_2_io_out_psum)
  );
  basic_PE PE_Array_0_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_3_clock),
    .reset(PE_Array_0_3_reset),
    .io_in_activate(PE_Array_0_3_io_in_activate),
    .io_in_weight(PE_Array_0_3_io_in_weight),
    .io_in_psum(PE_Array_0_3_io_in_psum),
    .io_in_flow(PE_Array_0_3_io_in_flow),
    .io_in_shift(PE_Array_0_3_io_in_shift),
    .io_out_activate(PE_Array_0_3_io_out_activate),
    .io_out_weight(PE_Array_0_3_io_out_weight),
    .io_out_psum(PE_Array_0_3_io_out_psum)
  );
  basic_PE PE_Array_0_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_4_clock),
    .reset(PE_Array_0_4_reset),
    .io_in_activate(PE_Array_0_4_io_in_activate),
    .io_in_weight(PE_Array_0_4_io_in_weight),
    .io_in_psum(PE_Array_0_4_io_in_psum),
    .io_in_flow(PE_Array_0_4_io_in_flow),
    .io_in_shift(PE_Array_0_4_io_in_shift),
    .io_out_activate(PE_Array_0_4_io_out_activate),
    .io_out_weight(PE_Array_0_4_io_out_weight),
    .io_out_psum(PE_Array_0_4_io_out_psum)
  );
  basic_PE PE_Array_0_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_5_clock),
    .reset(PE_Array_0_5_reset),
    .io_in_activate(PE_Array_0_5_io_in_activate),
    .io_in_weight(PE_Array_0_5_io_in_weight),
    .io_in_psum(PE_Array_0_5_io_in_psum),
    .io_in_flow(PE_Array_0_5_io_in_flow),
    .io_in_shift(PE_Array_0_5_io_in_shift),
    .io_out_activate(PE_Array_0_5_io_out_activate),
    .io_out_weight(PE_Array_0_5_io_out_weight),
    .io_out_psum(PE_Array_0_5_io_out_psum)
  );
  basic_PE PE_Array_0_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_6_clock),
    .reset(PE_Array_0_6_reset),
    .io_in_activate(PE_Array_0_6_io_in_activate),
    .io_in_weight(PE_Array_0_6_io_in_weight),
    .io_in_psum(PE_Array_0_6_io_in_psum),
    .io_in_flow(PE_Array_0_6_io_in_flow),
    .io_in_shift(PE_Array_0_6_io_in_shift),
    .io_out_activate(PE_Array_0_6_io_out_activate),
    .io_out_weight(PE_Array_0_6_io_out_weight),
    .io_out_psum(PE_Array_0_6_io_out_psum)
  );
  basic_PE PE_Array_0_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_7_clock),
    .reset(PE_Array_0_7_reset),
    .io_in_activate(PE_Array_0_7_io_in_activate),
    .io_in_weight(PE_Array_0_7_io_in_weight),
    .io_in_psum(PE_Array_0_7_io_in_psum),
    .io_in_flow(PE_Array_0_7_io_in_flow),
    .io_in_shift(PE_Array_0_7_io_in_shift),
    .io_out_activate(PE_Array_0_7_io_out_activate),
    .io_out_weight(PE_Array_0_7_io_out_weight),
    .io_out_psum(PE_Array_0_7_io_out_psum)
  );
  basic_PE PE_Array_0_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_8_clock),
    .reset(PE_Array_0_8_reset),
    .io_in_activate(PE_Array_0_8_io_in_activate),
    .io_in_weight(PE_Array_0_8_io_in_weight),
    .io_in_psum(PE_Array_0_8_io_in_psum),
    .io_in_flow(PE_Array_0_8_io_in_flow),
    .io_in_shift(PE_Array_0_8_io_in_shift),
    .io_out_activate(PE_Array_0_8_io_out_activate),
    .io_out_weight(PE_Array_0_8_io_out_weight),
    .io_out_psum(PE_Array_0_8_io_out_psum)
  );
  basic_PE PE_Array_0_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_9_clock),
    .reset(PE_Array_0_9_reset),
    .io_in_activate(PE_Array_0_9_io_in_activate),
    .io_in_weight(PE_Array_0_9_io_in_weight),
    .io_in_psum(PE_Array_0_9_io_in_psum),
    .io_in_flow(PE_Array_0_9_io_in_flow),
    .io_in_shift(PE_Array_0_9_io_in_shift),
    .io_out_activate(PE_Array_0_9_io_out_activate),
    .io_out_weight(PE_Array_0_9_io_out_weight),
    .io_out_psum(PE_Array_0_9_io_out_psum)
  );
  basic_PE PE_Array_0_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_10_clock),
    .reset(PE_Array_0_10_reset),
    .io_in_activate(PE_Array_0_10_io_in_activate),
    .io_in_weight(PE_Array_0_10_io_in_weight),
    .io_in_psum(PE_Array_0_10_io_in_psum),
    .io_in_flow(PE_Array_0_10_io_in_flow),
    .io_in_shift(PE_Array_0_10_io_in_shift),
    .io_out_activate(PE_Array_0_10_io_out_activate),
    .io_out_weight(PE_Array_0_10_io_out_weight),
    .io_out_psum(PE_Array_0_10_io_out_psum)
  );
  basic_PE PE_Array_0_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_11_clock),
    .reset(PE_Array_0_11_reset),
    .io_in_activate(PE_Array_0_11_io_in_activate),
    .io_in_weight(PE_Array_0_11_io_in_weight),
    .io_in_psum(PE_Array_0_11_io_in_psum),
    .io_in_flow(PE_Array_0_11_io_in_flow),
    .io_in_shift(PE_Array_0_11_io_in_shift),
    .io_out_activate(PE_Array_0_11_io_out_activate),
    .io_out_weight(PE_Array_0_11_io_out_weight),
    .io_out_psum(PE_Array_0_11_io_out_psum)
  );
  basic_PE PE_Array_0_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_12_clock),
    .reset(PE_Array_0_12_reset),
    .io_in_activate(PE_Array_0_12_io_in_activate),
    .io_in_weight(PE_Array_0_12_io_in_weight),
    .io_in_psum(PE_Array_0_12_io_in_psum),
    .io_in_flow(PE_Array_0_12_io_in_flow),
    .io_in_shift(PE_Array_0_12_io_in_shift),
    .io_out_activate(PE_Array_0_12_io_out_activate),
    .io_out_weight(PE_Array_0_12_io_out_weight),
    .io_out_psum(PE_Array_0_12_io_out_psum)
  );
  basic_PE PE_Array_0_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_13_clock),
    .reset(PE_Array_0_13_reset),
    .io_in_activate(PE_Array_0_13_io_in_activate),
    .io_in_weight(PE_Array_0_13_io_in_weight),
    .io_in_psum(PE_Array_0_13_io_in_psum),
    .io_in_flow(PE_Array_0_13_io_in_flow),
    .io_in_shift(PE_Array_0_13_io_in_shift),
    .io_out_activate(PE_Array_0_13_io_out_activate),
    .io_out_weight(PE_Array_0_13_io_out_weight),
    .io_out_psum(PE_Array_0_13_io_out_psum)
  );
  basic_PE PE_Array_0_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_14_clock),
    .reset(PE_Array_0_14_reset),
    .io_in_activate(PE_Array_0_14_io_in_activate),
    .io_in_weight(PE_Array_0_14_io_in_weight),
    .io_in_psum(PE_Array_0_14_io_in_psum),
    .io_in_flow(PE_Array_0_14_io_in_flow),
    .io_in_shift(PE_Array_0_14_io_in_shift),
    .io_out_activate(PE_Array_0_14_io_out_activate),
    .io_out_weight(PE_Array_0_14_io_out_weight),
    .io_out_psum(PE_Array_0_14_io_out_psum)
  );
  basic_PE PE_Array_0_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_15_clock),
    .reset(PE_Array_0_15_reset),
    .io_in_activate(PE_Array_0_15_io_in_activate),
    .io_in_weight(PE_Array_0_15_io_in_weight),
    .io_in_psum(PE_Array_0_15_io_in_psum),
    .io_in_flow(PE_Array_0_15_io_in_flow),
    .io_in_shift(PE_Array_0_15_io_in_shift),
    .io_out_activate(PE_Array_0_15_io_out_activate),
    .io_out_weight(PE_Array_0_15_io_out_weight),
    .io_out_psum(PE_Array_0_15_io_out_psum)
  );
  basic_PE PE_Array_0_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_16_clock),
    .reset(PE_Array_0_16_reset),
    .io_in_activate(PE_Array_0_16_io_in_activate),
    .io_in_weight(PE_Array_0_16_io_in_weight),
    .io_in_psum(PE_Array_0_16_io_in_psum),
    .io_in_flow(PE_Array_0_16_io_in_flow),
    .io_in_shift(PE_Array_0_16_io_in_shift),
    .io_out_activate(PE_Array_0_16_io_out_activate),
    .io_out_weight(PE_Array_0_16_io_out_weight),
    .io_out_psum(PE_Array_0_16_io_out_psum)
  );
  basic_PE PE_Array_0_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_17_clock),
    .reset(PE_Array_0_17_reset),
    .io_in_activate(PE_Array_0_17_io_in_activate),
    .io_in_weight(PE_Array_0_17_io_in_weight),
    .io_in_psum(PE_Array_0_17_io_in_psum),
    .io_in_flow(PE_Array_0_17_io_in_flow),
    .io_in_shift(PE_Array_0_17_io_in_shift),
    .io_out_activate(PE_Array_0_17_io_out_activate),
    .io_out_weight(PE_Array_0_17_io_out_weight),
    .io_out_psum(PE_Array_0_17_io_out_psum)
  );
  basic_PE PE_Array_0_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_18_clock),
    .reset(PE_Array_0_18_reset),
    .io_in_activate(PE_Array_0_18_io_in_activate),
    .io_in_weight(PE_Array_0_18_io_in_weight),
    .io_in_psum(PE_Array_0_18_io_in_psum),
    .io_in_flow(PE_Array_0_18_io_in_flow),
    .io_in_shift(PE_Array_0_18_io_in_shift),
    .io_out_activate(PE_Array_0_18_io_out_activate),
    .io_out_weight(PE_Array_0_18_io_out_weight),
    .io_out_psum(PE_Array_0_18_io_out_psum)
  );
  basic_PE PE_Array_0_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_19_clock),
    .reset(PE_Array_0_19_reset),
    .io_in_activate(PE_Array_0_19_io_in_activate),
    .io_in_weight(PE_Array_0_19_io_in_weight),
    .io_in_psum(PE_Array_0_19_io_in_psum),
    .io_in_flow(PE_Array_0_19_io_in_flow),
    .io_in_shift(PE_Array_0_19_io_in_shift),
    .io_out_activate(PE_Array_0_19_io_out_activate),
    .io_out_weight(PE_Array_0_19_io_out_weight),
    .io_out_psum(PE_Array_0_19_io_out_psum)
  );
  basic_PE PE_Array_0_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_20_clock),
    .reset(PE_Array_0_20_reset),
    .io_in_activate(PE_Array_0_20_io_in_activate),
    .io_in_weight(PE_Array_0_20_io_in_weight),
    .io_in_psum(PE_Array_0_20_io_in_psum),
    .io_in_flow(PE_Array_0_20_io_in_flow),
    .io_in_shift(PE_Array_0_20_io_in_shift),
    .io_out_activate(PE_Array_0_20_io_out_activate),
    .io_out_weight(PE_Array_0_20_io_out_weight),
    .io_out_psum(PE_Array_0_20_io_out_psum)
  );
  basic_PE PE_Array_0_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_21_clock),
    .reset(PE_Array_0_21_reset),
    .io_in_activate(PE_Array_0_21_io_in_activate),
    .io_in_weight(PE_Array_0_21_io_in_weight),
    .io_in_psum(PE_Array_0_21_io_in_psum),
    .io_in_flow(PE_Array_0_21_io_in_flow),
    .io_in_shift(PE_Array_0_21_io_in_shift),
    .io_out_activate(PE_Array_0_21_io_out_activate),
    .io_out_weight(PE_Array_0_21_io_out_weight),
    .io_out_psum(PE_Array_0_21_io_out_psum)
  );
  basic_PE PE_Array_0_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_22_clock),
    .reset(PE_Array_0_22_reset),
    .io_in_activate(PE_Array_0_22_io_in_activate),
    .io_in_weight(PE_Array_0_22_io_in_weight),
    .io_in_psum(PE_Array_0_22_io_in_psum),
    .io_in_flow(PE_Array_0_22_io_in_flow),
    .io_in_shift(PE_Array_0_22_io_in_shift),
    .io_out_activate(PE_Array_0_22_io_out_activate),
    .io_out_weight(PE_Array_0_22_io_out_weight),
    .io_out_psum(PE_Array_0_22_io_out_psum)
  );
  basic_PE PE_Array_0_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_23_clock),
    .reset(PE_Array_0_23_reset),
    .io_in_activate(PE_Array_0_23_io_in_activate),
    .io_in_weight(PE_Array_0_23_io_in_weight),
    .io_in_psum(PE_Array_0_23_io_in_psum),
    .io_in_flow(PE_Array_0_23_io_in_flow),
    .io_in_shift(PE_Array_0_23_io_in_shift),
    .io_out_activate(PE_Array_0_23_io_out_activate),
    .io_out_weight(PE_Array_0_23_io_out_weight),
    .io_out_psum(PE_Array_0_23_io_out_psum)
  );
  basic_PE PE_Array_0_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_24_clock),
    .reset(PE_Array_0_24_reset),
    .io_in_activate(PE_Array_0_24_io_in_activate),
    .io_in_weight(PE_Array_0_24_io_in_weight),
    .io_in_psum(PE_Array_0_24_io_in_psum),
    .io_in_flow(PE_Array_0_24_io_in_flow),
    .io_in_shift(PE_Array_0_24_io_in_shift),
    .io_out_activate(PE_Array_0_24_io_out_activate),
    .io_out_weight(PE_Array_0_24_io_out_weight),
    .io_out_psum(PE_Array_0_24_io_out_psum)
  );
  basic_PE PE_Array_0_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_25_clock),
    .reset(PE_Array_0_25_reset),
    .io_in_activate(PE_Array_0_25_io_in_activate),
    .io_in_weight(PE_Array_0_25_io_in_weight),
    .io_in_psum(PE_Array_0_25_io_in_psum),
    .io_in_flow(PE_Array_0_25_io_in_flow),
    .io_in_shift(PE_Array_0_25_io_in_shift),
    .io_out_activate(PE_Array_0_25_io_out_activate),
    .io_out_weight(PE_Array_0_25_io_out_weight),
    .io_out_psum(PE_Array_0_25_io_out_psum)
  );
  basic_PE PE_Array_0_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_26_clock),
    .reset(PE_Array_0_26_reset),
    .io_in_activate(PE_Array_0_26_io_in_activate),
    .io_in_weight(PE_Array_0_26_io_in_weight),
    .io_in_psum(PE_Array_0_26_io_in_psum),
    .io_in_flow(PE_Array_0_26_io_in_flow),
    .io_in_shift(PE_Array_0_26_io_in_shift),
    .io_out_activate(PE_Array_0_26_io_out_activate),
    .io_out_weight(PE_Array_0_26_io_out_weight),
    .io_out_psum(PE_Array_0_26_io_out_psum)
  );
  basic_PE PE_Array_0_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_27_clock),
    .reset(PE_Array_0_27_reset),
    .io_in_activate(PE_Array_0_27_io_in_activate),
    .io_in_weight(PE_Array_0_27_io_in_weight),
    .io_in_psum(PE_Array_0_27_io_in_psum),
    .io_in_flow(PE_Array_0_27_io_in_flow),
    .io_in_shift(PE_Array_0_27_io_in_shift),
    .io_out_activate(PE_Array_0_27_io_out_activate),
    .io_out_weight(PE_Array_0_27_io_out_weight),
    .io_out_psum(PE_Array_0_27_io_out_psum)
  );
  basic_PE PE_Array_0_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_28_clock),
    .reset(PE_Array_0_28_reset),
    .io_in_activate(PE_Array_0_28_io_in_activate),
    .io_in_weight(PE_Array_0_28_io_in_weight),
    .io_in_psum(PE_Array_0_28_io_in_psum),
    .io_in_flow(PE_Array_0_28_io_in_flow),
    .io_in_shift(PE_Array_0_28_io_in_shift),
    .io_out_activate(PE_Array_0_28_io_out_activate),
    .io_out_weight(PE_Array_0_28_io_out_weight),
    .io_out_psum(PE_Array_0_28_io_out_psum)
  );
  basic_PE PE_Array_0_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_29_clock),
    .reset(PE_Array_0_29_reset),
    .io_in_activate(PE_Array_0_29_io_in_activate),
    .io_in_weight(PE_Array_0_29_io_in_weight),
    .io_in_psum(PE_Array_0_29_io_in_psum),
    .io_in_flow(PE_Array_0_29_io_in_flow),
    .io_in_shift(PE_Array_0_29_io_in_shift),
    .io_out_activate(PE_Array_0_29_io_out_activate),
    .io_out_weight(PE_Array_0_29_io_out_weight),
    .io_out_psum(PE_Array_0_29_io_out_psum)
  );
  basic_PE PE_Array_0_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_30_clock),
    .reset(PE_Array_0_30_reset),
    .io_in_activate(PE_Array_0_30_io_in_activate),
    .io_in_weight(PE_Array_0_30_io_in_weight),
    .io_in_psum(PE_Array_0_30_io_in_psum),
    .io_in_flow(PE_Array_0_30_io_in_flow),
    .io_in_shift(PE_Array_0_30_io_in_shift),
    .io_out_activate(PE_Array_0_30_io_out_activate),
    .io_out_weight(PE_Array_0_30_io_out_weight),
    .io_out_psum(PE_Array_0_30_io_out_psum)
  );
  basic_PE PE_Array_0_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_31_clock),
    .reset(PE_Array_0_31_reset),
    .io_in_activate(PE_Array_0_31_io_in_activate),
    .io_in_weight(PE_Array_0_31_io_in_weight),
    .io_in_psum(PE_Array_0_31_io_in_psum),
    .io_in_flow(PE_Array_0_31_io_in_flow),
    .io_in_shift(PE_Array_0_31_io_in_shift),
    .io_out_activate(PE_Array_0_31_io_out_activate),
    .io_out_weight(PE_Array_0_31_io_out_weight),
    .io_out_psum(PE_Array_0_31_io_out_psum)
  );
  basic_PE PE_Array_1_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_0_clock),
    .reset(PE_Array_1_0_reset),
    .io_in_activate(PE_Array_1_0_io_in_activate),
    .io_in_weight(PE_Array_1_0_io_in_weight),
    .io_in_psum(PE_Array_1_0_io_in_psum),
    .io_in_flow(PE_Array_1_0_io_in_flow),
    .io_in_shift(PE_Array_1_0_io_in_shift),
    .io_out_activate(PE_Array_1_0_io_out_activate),
    .io_out_weight(PE_Array_1_0_io_out_weight),
    .io_out_psum(PE_Array_1_0_io_out_psum)
  );
  basic_PE PE_Array_1_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_1_clock),
    .reset(PE_Array_1_1_reset),
    .io_in_activate(PE_Array_1_1_io_in_activate),
    .io_in_weight(PE_Array_1_1_io_in_weight),
    .io_in_psum(PE_Array_1_1_io_in_psum),
    .io_in_flow(PE_Array_1_1_io_in_flow),
    .io_in_shift(PE_Array_1_1_io_in_shift),
    .io_out_activate(PE_Array_1_1_io_out_activate),
    .io_out_weight(PE_Array_1_1_io_out_weight),
    .io_out_psum(PE_Array_1_1_io_out_psum)
  );
  basic_PE PE_Array_1_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_2_clock),
    .reset(PE_Array_1_2_reset),
    .io_in_activate(PE_Array_1_2_io_in_activate),
    .io_in_weight(PE_Array_1_2_io_in_weight),
    .io_in_psum(PE_Array_1_2_io_in_psum),
    .io_in_flow(PE_Array_1_2_io_in_flow),
    .io_in_shift(PE_Array_1_2_io_in_shift),
    .io_out_activate(PE_Array_1_2_io_out_activate),
    .io_out_weight(PE_Array_1_2_io_out_weight),
    .io_out_psum(PE_Array_1_2_io_out_psum)
  );
  basic_PE PE_Array_1_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_3_clock),
    .reset(PE_Array_1_3_reset),
    .io_in_activate(PE_Array_1_3_io_in_activate),
    .io_in_weight(PE_Array_1_3_io_in_weight),
    .io_in_psum(PE_Array_1_3_io_in_psum),
    .io_in_flow(PE_Array_1_3_io_in_flow),
    .io_in_shift(PE_Array_1_3_io_in_shift),
    .io_out_activate(PE_Array_1_3_io_out_activate),
    .io_out_weight(PE_Array_1_3_io_out_weight),
    .io_out_psum(PE_Array_1_3_io_out_psum)
  );
  basic_PE PE_Array_1_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_4_clock),
    .reset(PE_Array_1_4_reset),
    .io_in_activate(PE_Array_1_4_io_in_activate),
    .io_in_weight(PE_Array_1_4_io_in_weight),
    .io_in_psum(PE_Array_1_4_io_in_psum),
    .io_in_flow(PE_Array_1_4_io_in_flow),
    .io_in_shift(PE_Array_1_4_io_in_shift),
    .io_out_activate(PE_Array_1_4_io_out_activate),
    .io_out_weight(PE_Array_1_4_io_out_weight),
    .io_out_psum(PE_Array_1_4_io_out_psum)
  );
  basic_PE PE_Array_1_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_5_clock),
    .reset(PE_Array_1_5_reset),
    .io_in_activate(PE_Array_1_5_io_in_activate),
    .io_in_weight(PE_Array_1_5_io_in_weight),
    .io_in_psum(PE_Array_1_5_io_in_psum),
    .io_in_flow(PE_Array_1_5_io_in_flow),
    .io_in_shift(PE_Array_1_5_io_in_shift),
    .io_out_activate(PE_Array_1_5_io_out_activate),
    .io_out_weight(PE_Array_1_5_io_out_weight),
    .io_out_psum(PE_Array_1_5_io_out_psum)
  );
  basic_PE PE_Array_1_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_6_clock),
    .reset(PE_Array_1_6_reset),
    .io_in_activate(PE_Array_1_6_io_in_activate),
    .io_in_weight(PE_Array_1_6_io_in_weight),
    .io_in_psum(PE_Array_1_6_io_in_psum),
    .io_in_flow(PE_Array_1_6_io_in_flow),
    .io_in_shift(PE_Array_1_6_io_in_shift),
    .io_out_activate(PE_Array_1_6_io_out_activate),
    .io_out_weight(PE_Array_1_6_io_out_weight),
    .io_out_psum(PE_Array_1_6_io_out_psum)
  );
  basic_PE PE_Array_1_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_7_clock),
    .reset(PE_Array_1_7_reset),
    .io_in_activate(PE_Array_1_7_io_in_activate),
    .io_in_weight(PE_Array_1_7_io_in_weight),
    .io_in_psum(PE_Array_1_7_io_in_psum),
    .io_in_flow(PE_Array_1_7_io_in_flow),
    .io_in_shift(PE_Array_1_7_io_in_shift),
    .io_out_activate(PE_Array_1_7_io_out_activate),
    .io_out_weight(PE_Array_1_7_io_out_weight),
    .io_out_psum(PE_Array_1_7_io_out_psum)
  );
  basic_PE PE_Array_1_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_8_clock),
    .reset(PE_Array_1_8_reset),
    .io_in_activate(PE_Array_1_8_io_in_activate),
    .io_in_weight(PE_Array_1_8_io_in_weight),
    .io_in_psum(PE_Array_1_8_io_in_psum),
    .io_in_flow(PE_Array_1_8_io_in_flow),
    .io_in_shift(PE_Array_1_8_io_in_shift),
    .io_out_activate(PE_Array_1_8_io_out_activate),
    .io_out_weight(PE_Array_1_8_io_out_weight),
    .io_out_psum(PE_Array_1_8_io_out_psum)
  );
  basic_PE PE_Array_1_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_9_clock),
    .reset(PE_Array_1_9_reset),
    .io_in_activate(PE_Array_1_9_io_in_activate),
    .io_in_weight(PE_Array_1_9_io_in_weight),
    .io_in_psum(PE_Array_1_9_io_in_psum),
    .io_in_flow(PE_Array_1_9_io_in_flow),
    .io_in_shift(PE_Array_1_9_io_in_shift),
    .io_out_activate(PE_Array_1_9_io_out_activate),
    .io_out_weight(PE_Array_1_9_io_out_weight),
    .io_out_psum(PE_Array_1_9_io_out_psum)
  );
  basic_PE PE_Array_1_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_10_clock),
    .reset(PE_Array_1_10_reset),
    .io_in_activate(PE_Array_1_10_io_in_activate),
    .io_in_weight(PE_Array_1_10_io_in_weight),
    .io_in_psum(PE_Array_1_10_io_in_psum),
    .io_in_flow(PE_Array_1_10_io_in_flow),
    .io_in_shift(PE_Array_1_10_io_in_shift),
    .io_out_activate(PE_Array_1_10_io_out_activate),
    .io_out_weight(PE_Array_1_10_io_out_weight),
    .io_out_psum(PE_Array_1_10_io_out_psum)
  );
  basic_PE PE_Array_1_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_11_clock),
    .reset(PE_Array_1_11_reset),
    .io_in_activate(PE_Array_1_11_io_in_activate),
    .io_in_weight(PE_Array_1_11_io_in_weight),
    .io_in_psum(PE_Array_1_11_io_in_psum),
    .io_in_flow(PE_Array_1_11_io_in_flow),
    .io_in_shift(PE_Array_1_11_io_in_shift),
    .io_out_activate(PE_Array_1_11_io_out_activate),
    .io_out_weight(PE_Array_1_11_io_out_weight),
    .io_out_psum(PE_Array_1_11_io_out_psum)
  );
  basic_PE PE_Array_1_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_12_clock),
    .reset(PE_Array_1_12_reset),
    .io_in_activate(PE_Array_1_12_io_in_activate),
    .io_in_weight(PE_Array_1_12_io_in_weight),
    .io_in_psum(PE_Array_1_12_io_in_psum),
    .io_in_flow(PE_Array_1_12_io_in_flow),
    .io_in_shift(PE_Array_1_12_io_in_shift),
    .io_out_activate(PE_Array_1_12_io_out_activate),
    .io_out_weight(PE_Array_1_12_io_out_weight),
    .io_out_psum(PE_Array_1_12_io_out_psum)
  );
  basic_PE PE_Array_1_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_13_clock),
    .reset(PE_Array_1_13_reset),
    .io_in_activate(PE_Array_1_13_io_in_activate),
    .io_in_weight(PE_Array_1_13_io_in_weight),
    .io_in_psum(PE_Array_1_13_io_in_psum),
    .io_in_flow(PE_Array_1_13_io_in_flow),
    .io_in_shift(PE_Array_1_13_io_in_shift),
    .io_out_activate(PE_Array_1_13_io_out_activate),
    .io_out_weight(PE_Array_1_13_io_out_weight),
    .io_out_psum(PE_Array_1_13_io_out_psum)
  );
  basic_PE PE_Array_1_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_14_clock),
    .reset(PE_Array_1_14_reset),
    .io_in_activate(PE_Array_1_14_io_in_activate),
    .io_in_weight(PE_Array_1_14_io_in_weight),
    .io_in_psum(PE_Array_1_14_io_in_psum),
    .io_in_flow(PE_Array_1_14_io_in_flow),
    .io_in_shift(PE_Array_1_14_io_in_shift),
    .io_out_activate(PE_Array_1_14_io_out_activate),
    .io_out_weight(PE_Array_1_14_io_out_weight),
    .io_out_psum(PE_Array_1_14_io_out_psum)
  );
  basic_PE PE_Array_1_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_15_clock),
    .reset(PE_Array_1_15_reset),
    .io_in_activate(PE_Array_1_15_io_in_activate),
    .io_in_weight(PE_Array_1_15_io_in_weight),
    .io_in_psum(PE_Array_1_15_io_in_psum),
    .io_in_flow(PE_Array_1_15_io_in_flow),
    .io_in_shift(PE_Array_1_15_io_in_shift),
    .io_out_activate(PE_Array_1_15_io_out_activate),
    .io_out_weight(PE_Array_1_15_io_out_weight),
    .io_out_psum(PE_Array_1_15_io_out_psum)
  );
  basic_PE PE_Array_1_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_16_clock),
    .reset(PE_Array_1_16_reset),
    .io_in_activate(PE_Array_1_16_io_in_activate),
    .io_in_weight(PE_Array_1_16_io_in_weight),
    .io_in_psum(PE_Array_1_16_io_in_psum),
    .io_in_flow(PE_Array_1_16_io_in_flow),
    .io_in_shift(PE_Array_1_16_io_in_shift),
    .io_out_activate(PE_Array_1_16_io_out_activate),
    .io_out_weight(PE_Array_1_16_io_out_weight),
    .io_out_psum(PE_Array_1_16_io_out_psum)
  );
  basic_PE PE_Array_1_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_17_clock),
    .reset(PE_Array_1_17_reset),
    .io_in_activate(PE_Array_1_17_io_in_activate),
    .io_in_weight(PE_Array_1_17_io_in_weight),
    .io_in_psum(PE_Array_1_17_io_in_psum),
    .io_in_flow(PE_Array_1_17_io_in_flow),
    .io_in_shift(PE_Array_1_17_io_in_shift),
    .io_out_activate(PE_Array_1_17_io_out_activate),
    .io_out_weight(PE_Array_1_17_io_out_weight),
    .io_out_psum(PE_Array_1_17_io_out_psum)
  );
  basic_PE PE_Array_1_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_18_clock),
    .reset(PE_Array_1_18_reset),
    .io_in_activate(PE_Array_1_18_io_in_activate),
    .io_in_weight(PE_Array_1_18_io_in_weight),
    .io_in_psum(PE_Array_1_18_io_in_psum),
    .io_in_flow(PE_Array_1_18_io_in_flow),
    .io_in_shift(PE_Array_1_18_io_in_shift),
    .io_out_activate(PE_Array_1_18_io_out_activate),
    .io_out_weight(PE_Array_1_18_io_out_weight),
    .io_out_psum(PE_Array_1_18_io_out_psum)
  );
  basic_PE PE_Array_1_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_19_clock),
    .reset(PE_Array_1_19_reset),
    .io_in_activate(PE_Array_1_19_io_in_activate),
    .io_in_weight(PE_Array_1_19_io_in_weight),
    .io_in_psum(PE_Array_1_19_io_in_psum),
    .io_in_flow(PE_Array_1_19_io_in_flow),
    .io_in_shift(PE_Array_1_19_io_in_shift),
    .io_out_activate(PE_Array_1_19_io_out_activate),
    .io_out_weight(PE_Array_1_19_io_out_weight),
    .io_out_psum(PE_Array_1_19_io_out_psum)
  );
  basic_PE PE_Array_1_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_20_clock),
    .reset(PE_Array_1_20_reset),
    .io_in_activate(PE_Array_1_20_io_in_activate),
    .io_in_weight(PE_Array_1_20_io_in_weight),
    .io_in_psum(PE_Array_1_20_io_in_psum),
    .io_in_flow(PE_Array_1_20_io_in_flow),
    .io_in_shift(PE_Array_1_20_io_in_shift),
    .io_out_activate(PE_Array_1_20_io_out_activate),
    .io_out_weight(PE_Array_1_20_io_out_weight),
    .io_out_psum(PE_Array_1_20_io_out_psum)
  );
  basic_PE PE_Array_1_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_21_clock),
    .reset(PE_Array_1_21_reset),
    .io_in_activate(PE_Array_1_21_io_in_activate),
    .io_in_weight(PE_Array_1_21_io_in_weight),
    .io_in_psum(PE_Array_1_21_io_in_psum),
    .io_in_flow(PE_Array_1_21_io_in_flow),
    .io_in_shift(PE_Array_1_21_io_in_shift),
    .io_out_activate(PE_Array_1_21_io_out_activate),
    .io_out_weight(PE_Array_1_21_io_out_weight),
    .io_out_psum(PE_Array_1_21_io_out_psum)
  );
  basic_PE PE_Array_1_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_22_clock),
    .reset(PE_Array_1_22_reset),
    .io_in_activate(PE_Array_1_22_io_in_activate),
    .io_in_weight(PE_Array_1_22_io_in_weight),
    .io_in_psum(PE_Array_1_22_io_in_psum),
    .io_in_flow(PE_Array_1_22_io_in_flow),
    .io_in_shift(PE_Array_1_22_io_in_shift),
    .io_out_activate(PE_Array_1_22_io_out_activate),
    .io_out_weight(PE_Array_1_22_io_out_weight),
    .io_out_psum(PE_Array_1_22_io_out_psum)
  );
  basic_PE PE_Array_1_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_23_clock),
    .reset(PE_Array_1_23_reset),
    .io_in_activate(PE_Array_1_23_io_in_activate),
    .io_in_weight(PE_Array_1_23_io_in_weight),
    .io_in_psum(PE_Array_1_23_io_in_psum),
    .io_in_flow(PE_Array_1_23_io_in_flow),
    .io_in_shift(PE_Array_1_23_io_in_shift),
    .io_out_activate(PE_Array_1_23_io_out_activate),
    .io_out_weight(PE_Array_1_23_io_out_weight),
    .io_out_psum(PE_Array_1_23_io_out_psum)
  );
  basic_PE PE_Array_1_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_24_clock),
    .reset(PE_Array_1_24_reset),
    .io_in_activate(PE_Array_1_24_io_in_activate),
    .io_in_weight(PE_Array_1_24_io_in_weight),
    .io_in_psum(PE_Array_1_24_io_in_psum),
    .io_in_flow(PE_Array_1_24_io_in_flow),
    .io_in_shift(PE_Array_1_24_io_in_shift),
    .io_out_activate(PE_Array_1_24_io_out_activate),
    .io_out_weight(PE_Array_1_24_io_out_weight),
    .io_out_psum(PE_Array_1_24_io_out_psum)
  );
  basic_PE PE_Array_1_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_25_clock),
    .reset(PE_Array_1_25_reset),
    .io_in_activate(PE_Array_1_25_io_in_activate),
    .io_in_weight(PE_Array_1_25_io_in_weight),
    .io_in_psum(PE_Array_1_25_io_in_psum),
    .io_in_flow(PE_Array_1_25_io_in_flow),
    .io_in_shift(PE_Array_1_25_io_in_shift),
    .io_out_activate(PE_Array_1_25_io_out_activate),
    .io_out_weight(PE_Array_1_25_io_out_weight),
    .io_out_psum(PE_Array_1_25_io_out_psum)
  );
  basic_PE PE_Array_1_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_26_clock),
    .reset(PE_Array_1_26_reset),
    .io_in_activate(PE_Array_1_26_io_in_activate),
    .io_in_weight(PE_Array_1_26_io_in_weight),
    .io_in_psum(PE_Array_1_26_io_in_psum),
    .io_in_flow(PE_Array_1_26_io_in_flow),
    .io_in_shift(PE_Array_1_26_io_in_shift),
    .io_out_activate(PE_Array_1_26_io_out_activate),
    .io_out_weight(PE_Array_1_26_io_out_weight),
    .io_out_psum(PE_Array_1_26_io_out_psum)
  );
  basic_PE PE_Array_1_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_27_clock),
    .reset(PE_Array_1_27_reset),
    .io_in_activate(PE_Array_1_27_io_in_activate),
    .io_in_weight(PE_Array_1_27_io_in_weight),
    .io_in_psum(PE_Array_1_27_io_in_psum),
    .io_in_flow(PE_Array_1_27_io_in_flow),
    .io_in_shift(PE_Array_1_27_io_in_shift),
    .io_out_activate(PE_Array_1_27_io_out_activate),
    .io_out_weight(PE_Array_1_27_io_out_weight),
    .io_out_psum(PE_Array_1_27_io_out_psum)
  );
  basic_PE PE_Array_1_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_28_clock),
    .reset(PE_Array_1_28_reset),
    .io_in_activate(PE_Array_1_28_io_in_activate),
    .io_in_weight(PE_Array_1_28_io_in_weight),
    .io_in_psum(PE_Array_1_28_io_in_psum),
    .io_in_flow(PE_Array_1_28_io_in_flow),
    .io_in_shift(PE_Array_1_28_io_in_shift),
    .io_out_activate(PE_Array_1_28_io_out_activate),
    .io_out_weight(PE_Array_1_28_io_out_weight),
    .io_out_psum(PE_Array_1_28_io_out_psum)
  );
  basic_PE PE_Array_1_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_29_clock),
    .reset(PE_Array_1_29_reset),
    .io_in_activate(PE_Array_1_29_io_in_activate),
    .io_in_weight(PE_Array_1_29_io_in_weight),
    .io_in_psum(PE_Array_1_29_io_in_psum),
    .io_in_flow(PE_Array_1_29_io_in_flow),
    .io_in_shift(PE_Array_1_29_io_in_shift),
    .io_out_activate(PE_Array_1_29_io_out_activate),
    .io_out_weight(PE_Array_1_29_io_out_weight),
    .io_out_psum(PE_Array_1_29_io_out_psum)
  );
  basic_PE PE_Array_1_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_30_clock),
    .reset(PE_Array_1_30_reset),
    .io_in_activate(PE_Array_1_30_io_in_activate),
    .io_in_weight(PE_Array_1_30_io_in_weight),
    .io_in_psum(PE_Array_1_30_io_in_psum),
    .io_in_flow(PE_Array_1_30_io_in_flow),
    .io_in_shift(PE_Array_1_30_io_in_shift),
    .io_out_activate(PE_Array_1_30_io_out_activate),
    .io_out_weight(PE_Array_1_30_io_out_weight),
    .io_out_psum(PE_Array_1_30_io_out_psum)
  );
  basic_PE PE_Array_1_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_31_clock),
    .reset(PE_Array_1_31_reset),
    .io_in_activate(PE_Array_1_31_io_in_activate),
    .io_in_weight(PE_Array_1_31_io_in_weight),
    .io_in_psum(PE_Array_1_31_io_in_psum),
    .io_in_flow(PE_Array_1_31_io_in_flow),
    .io_in_shift(PE_Array_1_31_io_in_shift),
    .io_out_activate(PE_Array_1_31_io_out_activate),
    .io_out_weight(PE_Array_1_31_io_out_weight),
    .io_out_psum(PE_Array_1_31_io_out_psum)
  );
  basic_PE PE_Array_2_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_0_clock),
    .reset(PE_Array_2_0_reset),
    .io_in_activate(PE_Array_2_0_io_in_activate),
    .io_in_weight(PE_Array_2_0_io_in_weight),
    .io_in_psum(PE_Array_2_0_io_in_psum),
    .io_in_flow(PE_Array_2_0_io_in_flow),
    .io_in_shift(PE_Array_2_0_io_in_shift),
    .io_out_activate(PE_Array_2_0_io_out_activate),
    .io_out_weight(PE_Array_2_0_io_out_weight),
    .io_out_psum(PE_Array_2_0_io_out_psum)
  );
  basic_PE PE_Array_2_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_1_clock),
    .reset(PE_Array_2_1_reset),
    .io_in_activate(PE_Array_2_1_io_in_activate),
    .io_in_weight(PE_Array_2_1_io_in_weight),
    .io_in_psum(PE_Array_2_1_io_in_psum),
    .io_in_flow(PE_Array_2_1_io_in_flow),
    .io_in_shift(PE_Array_2_1_io_in_shift),
    .io_out_activate(PE_Array_2_1_io_out_activate),
    .io_out_weight(PE_Array_2_1_io_out_weight),
    .io_out_psum(PE_Array_2_1_io_out_psum)
  );
  basic_PE PE_Array_2_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_2_clock),
    .reset(PE_Array_2_2_reset),
    .io_in_activate(PE_Array_2_2_io_in_activate),
    .io_in_weight(PE_Array_2_2_io_in_weight),
    .io_in_psum(PE_Array_2_2_io_in_psum),
    .io_in_flow(PE_Array_2_2_io_in_flow),
    .io_in_shift(PE_Array_2_2_io_in_shift),
    .io_out_activate(PE_Array_2_2_io_out_activate),
    .io_out_weight(PE_Array_2_2_io_out_weight),
    .io_out_psum(PE_Array_2_2_io_out_psum)
  );
  basic_PE PE_Array_2_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_3_clock),
    .reset(PE_Array_2_3_reset),
    .io_in_activate(PE_Array_2_3_io_in_activate),
    .io_in_weight(PE_Array_2_3_io_in_weight),
    .io_in_psum(PE_Array_2_3_io_in_psum),
    .io_in_flow(PE_Array_2_3_io_in_flow),
    .io_in_shift(PE_Array_2_3_io_in_shift),
    .io_out_activate(PE_Array_2_3_io_out_activate),
    .io_out_weight(PE_Array_2_3_io_out_weight),
    .io_out_psum(PE_Array_2_3_io_out_psum)
  );
  basic_PE PE_Array_2_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_4_clock),
    .reset(PE_Array_2_4_reset),
    .io_in_activate(PE_Array_2_4_io_in_activate),
    .io_in_weight(PE_Array_2_4_io_in_weight),
    .io_in_psum(PE_Array_2_4_io_in_psum),
    .io_in_flow(PE_Array_2_4_io_in_flow),
    .io_in_shift(PE_Array_2_4_io_in_shift),
    .io_out_activate(PE_Array_2_4_io_out_activate),
    .io_out_weight(PE_Array_2_4_io_out_weight),
    .io_out_psum(PE_Array_2_4_io_out_psum)
  );
  basic_PE PE_Array_2_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_5_clock),
    .reset(PE_Array_2_5_reset),
    .io_in_activate(PE_Array_2_5_io_in_activate),
    .io_in_weight(PE_Array_2_5_io_in_weight),
    .io_in_psum(PE_Array_2_5_io_in_psum),
    .io_in_flow(PE_Array_2_5_io_in_flow),
    .io_in_shift(PE_Array_2_5_io_in_shift),
    .io_out_activate(PE_Array_2_5_io_out_activate),
    .io_out_weight(PE_Array_2_5_io_out_weight),
    .io_out_psum(PE_Array_2_5_io_out_psum)
  );
  basic_PE PE_Array_2_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_6_clock),
    .reset(PE_Array_2_6_reset),
    .io_in_activate(PE_Array_2_6_io_in_activate),
    .io_in_weight(PE_Array_2_6_io_in_weight),
    .io_in_psum(PE_Array_2_6_io_in_psum),
    .io_in_flow(PE_Array_2_6_io_in_flow),
    .io_in_shift(PE_Array_2_6_io_in_shift),
    .io_out_activate(PE_Array_2_6_io_out_activate),
    .io_out_weight(PE_Array_2_6_io_out_weight),
    .io_out_psum(PE_Array_2_6_io_out_psum)
  );
  basic_PE PE_Array_2_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_7_clock),
    .reset(PE_Array_2_7_reset),
    .io_in_activate(PE_Array_2_7_io_in_activate),
    .io_in_weight(PE_Array_2_7_io_in_weight),
    .io_in_psum(PE_Array_2_7_io_in_psum),
    .io_in_flow(PE_Array_2_7_io_in_flow),
    .io_in_shift(PE_Array_2_7_io_in_shift),
    .io_out_activate(PE_Array_2_7_io_out_activate),
    .io_out_weight(PE_Array_2_7_io_out_weight),
    .io_out_psum(PE_Array_2_7_io_out_psum)
  );
  basic_PE PE_Array_2_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_8_clock),
    .reset(PE_Array_2_8_reset),
    .io_in_activate(PE_Array_2_8_io_in_activate),
    .io_in_weight(PE_Array_2_8_io_in_weight),
    .io_in_psum(PE_Array_2_8_io_in_psum),
    .io_in_flow(PE_Array_2_8_io_in_flow),
    .io_in_shift(PE_Array_2_8_io_in_shift),
    .io_out_activate(PE_Array_2_8_io_out_activate),
    .io_out_weight(PE_Array_2_8_io_out_weight),
    .io_out_psum(PE_Array_2_8_io_out_psum)
  );
  basic_PE PE_Array_2_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_9_clock),
    .reset(PE_Array_2_9_reset),
    .io_in_activate(PE_Array_2_9_io_in_activate),
    .io_in_weight(PE_Array_2_9_io_in_weight),
    .io_in_psum(PE_Array_2_9_io_in_psum),
    .io_in_flow(PE_Array_2_9_io_in_flow),
    .io_in_shift(PE_Array_2_9_io_in_shift),
    .io_out_activate(PE_Array_2_9_io_out_activate),
    .io_out_weight(PE_Array_2_9_io_out_weight),
    .io_out_psum(PE_Array_2_9_io_out_psum)
  );
  basic_PE PE_Array_2_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_10_clock),
    .reset(PE_Array_2_10_reset),
    .io_in_activate(PE_Array_2_10_io_in_activate),
    .io_in_weight(PE_Array_2_10_io_in_weight),
    .io_in_psum(PE_Array_2_10_io_in_psum),
    .io_in_flow(PE_Array_2_10_io_in_flow),
    .io_in_shift(PE_Array_2_10_io_in_shift),
    .io_out_activate(PE_Array_2_10_io_out_activate),
    .io_out_weight(PE_Array_2_10_io_out_weight),
    .io_out_psum(PE_Array_2_10_io_out_psum)
  );
  basic_PE PE_Array_2_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_11_clock),
    .reset(PE_Array_2_11_reset),
    .io_in_activate(PE_Array_2_11_io_in_activate),
    .io_in_weight(PE_Array_2_11_io_in_weight),
    .io_in_psum(PE_Array_2_11_io_in_psum),
    .io_in_flow(PE_Array_2_11_io_in_flow),
    .io_in_shift(PE_Array_2_11_io_in_shift),
    .io_out_activate(PE_Array_2_11_io_out_activate),
    .io_out_weight(PE_Array_2_11_io_out_weight),
    .io_out_psum(PE_Array_2_11_io_out_psum)
  );
  basic_PE PE_Array_2_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_12_clock),
    .reset(PE_Array_2_12_reset),
    .io_in_activate(PE_Array_2_12_io_in_activate),
    .io_in_weight(PE_Array_2_12_io_in_weight),
    .io_in_psum(PE_Array_2_12_io_in_psum),
    .io_in_flow(PE_Array_2_12_io_in_flow),
    .io_in_shift(PE_Array_2_12_io_in_shift),
    .io_out_activate(PE_Array_2_12_io_out_activate),
    .io_out_weight(PE_Array_2_12_io_out_weight),
    .io_out_psum(PE_Array_2_12_io_out_psum)
  );
  basic_PE PE_Array_2_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_13_clock),
    .reset(PE_Array_2_13_reset),
    .io_in_activate(PE_Array_2_13_io_in_activate),
    .io_in_weight(PE_Array_2_13_io_in_weight),
    .io_in_psum(PE_Array_2_13_io_in_psum),
    .io_in_flow(PE_Array_2_13_io_in_flow),
    .io_in_shift(PE_Array_2_13_io_in_shift),
    .io_out_activate(PE_Array_2_13_io_out_activate),
    .io_out_weight(PE_Array_2_13_io_out_weight),
    .io_out_psum(PE_Array_2_13_io_out_psum)
  );
  basic_PE PE_Array_2_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_14_clock),
    .reset(PE_Array_2_14_reset),
    .io_in_activate(PE_Array_2_14_io_in_activate),
    .io_in_weight(PE_Array_2_14_io_in_weight),
    .io_in_psum(PE_Array_2_14_io_in_psum),
    .io_in_flow(PE_Array_2_14_io_in_flow),
    .io_in_shift(PE_Array_2_14_io_in_shift),
    .io_out_activate(PE_Array_2_14_io_out_activate),
    .io_out_weight(PE_Array_2_14_io_out_weight),
    .io_out_psum(PE_Array_2_14_io_out_psum)
  );
  basic_PE PE_Array_2_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_15_clock),
    .reset(PE_Array_2_15_reset),
    .io_in_activate(PE_Array_2_15_io_in_activate),
    .io_in_weight(PE_Array_2_15_io_in_weight),
    .io_in_psum(PE_Array_2_15_io_in_psum),
    .io_in_flow(PE_Array_2_15_io_in_flow),
    .io_in_shift(PE_Array_2_15_io_in_shift),
    .io_out_activate(PE_Array_2_15_io_out_activate),
    .io_out_weight(PE_Array_2_15_io_out_weight),
    .io_out_psum(PE_Array_2_15_io_out_psum)
  );
  basic_PE PE_Array_2_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_16_clock),
    .reset(PE_Array_2_16_reset),
    .io_in_activate(PE_Array_2_16_io_in_activate),
    .io_in_weight(PE_Array_2_16_io_in_weight),
    .io_in_psum(PE_Array_2_16_io_in_psum),
    .io_in_flow(PE_Array_2_16_io_in_flow),
    .io_in_shift(PE_Array_2_16_io_in_shift),
    .io_out_activate(PE_Array_2_16_io_out_activate),
    .io_out_weight(PE_Array_2_16_io_out_weight),
    .io_out_psum(PE_Array_2_16_io_out_psum)
  );
  basic_PE PE_Array_2_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_17_clock),
    .reset(PE_Array_2_17_reset),
    .io_in_activate(PE_Array_2_17_io_in_activate),
    .io_in_weight(PE_Array_2_17_io_in_weight),
    .io_in_psum(PE_Array_2_17_io_in_psum),
    .io_in_flow(PE_Array_2_17_io_in_flow),
    .io_in_shift(PE_Array_2_17_io_in_shift),
    .io_out_activate(PE_Array_2_17_io_out_activate),
    .io_out_weight(PE_Array_2_17_io_out_weight),
    .io_out_psum(PE_Array_2_17_io_out_psum)
  );
  basic_PE PE_Array_2_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_18_clock),
    .reset(PE_Array_2_18_reset),
    .io_in_activate(PE_Array_2_18_io_in_activate),
    .io_in_weight(PE_Array_2_18_io_in_weight),
    .io_in_psum(PE_Array_2_18_io_in_psum),
    .io_in_flow(PE_Array_2_18_io_in_flow),
    .io_in_shift(PE_Array_2_18_io_in_shift),
    .io_out_activate(PE_Array_2_18_io_out_activate),
    .io_out_weight(PE_Array_2_18_io_out_weight),
    .io_out_psum(PE_Array_2_18_io_out_psum)
  );
  basic_PE PE_Array_2_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_19_clock),
    .reset(PE_Array_2_19_reset),
    .io_in_activate(PE_Array_2_19_io_in_activate),
    .io_in_weight(PE_Array_2_19_io_in_weight),
    .io_in_psum(PE_Array_2_19_io_in_psum),
    .io_in_flow(PE_Array_2_19_io_in_flow),
    .io_in_shift(PE_Array_2_19_io_in_shift),
    .io_out_activate(PE_Array_2_19_io_out_activate),
    .io_out_weight(PE_Array_2_19_io_out_weight),
    .io_out_psum(PE_Array_2_19_io_out_psum)
  );
  basic_PE PE_Array_2_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_20_clock),
    .reset(PE_Array_2_20_reset),
    .io_in_activate(PE_Array_2_20_io_in_activate),
    .io_in_weight(PE_Array_2_20_io_in_weight),
    .io_in_psum(PE_Array_2_20_io_in_psum),
    .io_in_flow(PE_Array_2_20_io_in_flow),
    .io_in_shift(PE_Array_2_20_io_in_shift),
    .io_out_activate(PE_Array_2_20_io_out_activate),
    .io_out_weight(PE_Array_2_20_io_out_weight),
    .io_out_psum(PE_Array_2_20_io_out_psum)
  );
  basic_PE PE_Array_2_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_21_clock),
    .reset(PE_Array_2_21_reset),
    .io_in_activate(PE_Array_2_21_io_in_activate),
    .io_in_weight(PE_Array_2_21_io_in_weight),
    .io_in_psum(PE_Array_2_21_io_in_psum),
    .io_in_flow(PE_Array_2_21_io_in_flow),
    .io_in_shift(PE_Array_2_21_io_in_shift),
    .io_out_activate(PE_Array_2_21_io_out_activate),
    .io_out_weight(PE_Array_2_21_io_out_weight),
    .io_out_psum(PE_Array_2_21_io_out_psum)
  );
  basic_PE PE_Array_2_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_22_clock),
    .reset(PE_Array_2_22_reset),
    .io_in_activate(PE_Array_2_22_io_in_activate),
    .io_in_weight(PE_Array_2_22_io_in_weight),
    .io_in_psum(PE_Array_2_22_io_in_psum),
    .io_in_flow(PE_Array_2_22_io_in_flow),
    .io_in_shift(PE_Array_2_22_io_in_shift),
    .io_out_activate(PE_Array_2_22_io_out_activate),
    .io_out_weight(PE_Array_2_22_io_out_weight),
    .io_out_psum(PE_Array_2_22_io_out_psum)
  );
  basic_PE PE_Array_2_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_23_clock),
    .reset(PE_Array_2_23_reset),
    .io_in_activate(PE_Array_2_23_io_in_activate),
    .io_in_weight(PE_Array_2_23_io_in_weight),
    .io_in_psum(PE_Array_2_23_io_in_psum),
    .io_in_flow(PE_Array_2_23_io_in_flow),
    .io_in_shift(PE_Array_2_23_io_in_shift),
    .io_out_activate(PE_Array_2_23_io_out_activate),
    .io_out_weight(PE_Array_2_23_io_out_weight),
    .io_out_psum(PE_Array_2_23_io_out_psum)
  );
  basic_PE PE_Array_2_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_24_clock),
    .reset(PE_Array_2_24_reset),
    .io_in_activate(PE_Array_2_24_io_in_activate),
    .io_in_weight(PE_Array_2_24_io_in_weight),
    .io_in_psum(PE_Array_2_24_io_in_psum),
    .io_in_flow(PE_Array_2_24_io_in_flow),
    .io_in_shift(PE_Array_2_24_io_in_shift),
    .io_out_activate(PE_Array_2_24_io_out_activate),
    .io_out_weight(PE_Array_2_24_io_out_weight),
    .io_out_psum(PE_Array_2_24_io_out_psum)
  );
  basic_PE PE_Array_2_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_25_clock),
    .reset(PE_Array_2_25_reset),
    .io_in_activate(PE_Array_2_25_io_in_activate),
    .io_in_weight(PE_Array_2_25_io_in_weight),
    .io_in_psum(PE_Array_2_25_io_in_psum),
    .io_in_flow(PE_Array_2_25_io_in_flow),
    .io_in_shift(PE_Array_2_25_io_in_shift),
    .io_out_activate(PE_Array_2_25_io_out_activate),
    .io_out_weight(PE_Array_2_25_io_out_weight),
    .io_out_psum(PE_Array_2_25_io_out_psum)
  );
  basic_PE PE_Array_2_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_26_clock),
    .reset(PE_Array_2_26_reset),
    .io_in_activate(PE_Array_2_26_io_in_activate),
    .io_in_weight(PE_Array_2_26_io_in_weight),
    .io_in_psum(PE_Array_2_26_io_in_psum),
    .io_in_flow(PE_Array_2_26_io_in_flow),
    .io_in_shift(PE_Array_2_26_io_in_shift),
    .io_out_activate(PE_Array_2_26_io_out_activate),
    .io_out_weight(PE_Array_2_26_io_out_weight),
    .io_out_psum(PE_Array_2_26_io_out_psum)
  );
  basic_PE PE_Array_2_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_27_clock),
    .reset(PE_Array_2_27_reset),
    .io_in_activate(PE_Array_2_27_io_in_activate),
    .io_in_weight(PE_Array_2_27_io_in_weight),
    .io_in_psum(PE_Array_2_27_io_in_psum),
    .io_in_flow(PE_Array_2_27_io_in_flow),
    .io_in_shift(PE_Array_2_27_io_in_shift),
    .io_out_activate(PE_Array_2_27_io_out_activate),
    .io_out_weight(PE_Array_2_27_io_out_weight),
    .io_out_psum(PE_Array_2_27_io_out_psum)
  );
  basic_PE PE_Array_2_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_28_clock),
    .reset(PE_Array_2_28_reset),
    .io_in_activate(PE_Array_2_28_io_in_activate),
    .io_in_weight(PE_Array_2_28_io_in_weight),
    .io_in_psum(PE_Array_2_28_io_in_psum),
    .io_in_flow(PE_Array_2_28_io_in_flow),
    .io_in_shift(PE_Array_2_28_io_in_shift),
    .io_out_activate(PE_Array_2_28_io_out_activate),
    .io_out_weight(PE_Array_2_28_io_out_weight),
    .io_out_psum(PE_Array_2_28_io_out_psum)
  );
  basic_PE PE_Array_2_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_29_clock),
    .reset(PE_Array_2_29_reset),
    .io_in_activate(PE_Array_2_29_io_in_activate),
    .io_in_weight(PE_Array_2_29_io_in_weight),
    .io_in_psum(PE_Array_2_29_io_in_psum),
    .io_in_flow(PE_Array_2_29_io_in_flow),
    .io_in_shift(PE_Array_2_29_io_in_shift),
    .io_out_activate(PE_Array_2_29_io_out_activate),
    .io_out_weight(PE_Array_2_29_io_out_weight),
    .io_out_psum(PE_Array_2_29_io_out_psum)
  );
  basic_PE PE_Array_2_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_30_clock),
    .reset(PE_Array_2_30_reset),
    .io_in_activate(PE_Array_2_30_io_in_activate),
    .io_in_weight(PE_Array_2_30_io_in_weight),
    .io_in_psum(PE_Array_2_30_io_in_psum),
    .io_in_flow(PE_Array_2_30_io_in_flow),
    .io_in_shift(PE_Array_2_30_io_in_shift),
    .io_out_activate(PE_Array_2_30_io_out_activate),
    .io_out_weight(PE_Array_2_30_io_out_weight),
    .io_out_psum(PE_Array_2_30_io_out_psum)
  );
  basic_PE PE_Array_2_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_31_clock),
    .reset(PE_Array_2_31_reset),
    .io_in_activate(PE_Array_2_31_io_in_activate),
    .io_in_weight(PE_Array_2_31_io_in_weight),
    .io_in_psum(PE_Array_2_31_io_in_psum),
    .io_in_flow(PE_Array_2_31_io_in_flow),
    .io_in_shift(PE_Array_2_31_io_in_shift),
    .io_out_activate(PE_Array_2_31_io_out_activate),
    .io_out_weight(PE_Array_2_31_io_out_weight),
    .io_out_psum(PE_Array_2_31_io_out_psum)
  );
  basic_PE PE_Array_3_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_0_clock),
    .reset(PE_Array_3_0_reset),
    .io_in_activate(PE_Array_3_0_io_in_activate),
    .io_in_weight(PE_Array_3_0_io_in_weight),
    .io_in_psum(PE_Array_3_0_io_in_psum),
    .io_in_flow(PE_Array_3_0_io_in_flow),
    .io_in_shift(PE_Array_3_0_io_in_shift),
    .io_out_activate(PE_Array_3_0_io_out_activate),
    .io_out_weight(PE_Array_3_0_io_out_weight),
    .io_out_psum(PE_Array_3_0_io_out_psum)
  );
  basic_PE PE_Array_3_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_1_clock),
    .reset(PE_Array_3_1_reset),
    .io_in_activate(PE_Array_3_1_io_in_activate),
    .io_in_weight(PE_Array_3_1_io_in_weight),
    .io_in_psum(PE_Array_3_1_io_in_psum),
    .io_in_flow(PE_Array_3_1_io_in_flow),
    .io_in_shift(PE_Array_3_1_io_in_shift),
    .io_out_activate(PE_Array_3_1_io_out_activate),
    .io_out_weight(PE_Array_3_1_io_out_weight),
    .io_out_psum(PE_Array_3_1_io_out_psum)
  );
  basic_PE PE_Array_3_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_2_clock),
    .reset(PE_Array_3_2_reset),
    .io_in_activate(PE_Array_3_2_io_in_activate),
    .io_in_weight(PE_Array_3_2_io_in_weight),
    .io_in_psum(PE_Array_3_2_io_in_psum),
    .io_in_flow(PE_Array_3_2_io_in_flow),
    .io_in_shift(PE_Array_3_2_io_in_shift),
    .io_out_activate(PE_Array_3_2_io_out_activate),
    .io_out_weight(PE_Array_3_2_io_out_weight),
    .io_out_psum(PE_Array_3_2_io_out_psum)
  );
  basic_PE PE_Array_3_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_3_clock),
    .reset(PE_Array_3_3_reset),
    .io_in_activate(PE_Array_3_3_io_in_activate),
    .io_in_weight(PE_Array_3_3_io_in_weight),
    .io_in_psum(PE_Array_3_3_io_in_psum),
    .io_in_flow(PE_Array_3_3_io_in_flow),
    .io_in_shift(PE_Array_3_3_io_in_shift),
    .io_out_activate(PE_Array_3_3_io_out_activate),
    .io_out_weight(PE_Array_3_3_io_out_weight),
    .io_out_psum(PE_Array_3_3_io_out_psum)
  );
  basic_PE PE_Array_3_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_4_clock),
    .reset(PE_Array_3_4_reset),
    .io_in_activate(PE_Array_3_4_io_in_activate),
    .io_in_weight(PE_Array_3_4_io_in_weight),
    .io_in_psum(PE_Array_3_4_io_in_psum),
    .io_in_flow(PE_Array_3_4_io_in_flow),
    .io_in_shift(PE_Array_3_4_io_in_shift),
    .io_out_activate(PE_Array_3_4_io_out_activate),
    .io_out_weight(PE_Array_3_4_io_out_weight),
    .io_out_psum(PE_Array_3_4_io_out_psum)
  );
  basic_PE PE_Array_3_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_5_clock),
    .reset(PE_Array_3_5_reset),
    .io_in_activate(PE_Array_3_5_io_in_activate),
    .io_in_weight(PE_Array_3_5_io_in_weight),
    .io_in_psum(PE_Array_3_5_io_in_psum),
    .io_in_flow(PE_Array_3_5_io_in_flow),
    .io_in_shift(PE_Array_3_5_io_in_shift),
    .io_out_activate(PE_Array_3_5_io_out_activate),
    .io_out_weight(PE_Array_3_5_io_out_weight),
    .io_out_psum(PE_Array_3_5_io_out_psum)
  );
  basic_PE PE_Array_3_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_6_clock),
    .reset(PE_Array_3_6_reset),
    .io_in_activate(PE_Array_3_6_io_in_activate),
    .io_in_weight(PE_Array_3_6_io_in_weight),
    .io_in_psum(PE_Array_3_6_io_in_psum),
    .io_in_flow(PE_Array_3_6_io_in_flow),
    .io_in_shift(PE_Array_3_6_io_in_shift),
    .io_out_activate(PE_Array_3_6_io_out_activate),
    .io_out_weight(PE_Array_3_6_io_out_weight),
    .io_out_psum(PE_Array_3_6_io_out_psum)
  );
  basic_PE PE_Array_3_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_7_clock),
    .reset(PE_Array_3_7_reset),
    .io_in_activate(PE_Array_3_7_io_in_activate),
    .io_in_weight(PE_Array_3_7_io_in_weight),
    .io_in_psum(PE_Array_3_7_io_in_psum),
    .io_in_flow(PE_Array_3_7_io_in_flow),
    .io_in_shift(PE_Array_3_7_io_in_shift),
    .io_out_activate(PE_Array_3_7_io_out_activate),
    .io_out_weight(PE_Array_3_7_io_out_weight),
    .io_out_psum(PE_Array_3_7_io_out_psum)
  );
  basic_PE PE_Array_3_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_8_clock),
    .reset(PE_Array_3_8_reset),
    .io_in_activate(PE_Array_3_8_io_in_activate),
    .io_in_weight(PE_Array_3_8_io_in_weight),
    .io_in_psum(PE_Array_3_8_io_in_psum),
    .io_in_flow(PE_Array_3_8_io_in_flow),
    .io_in_shift(PE_Array_3_8_io_in_shift),
    .io_out_activate(PE_Array_3_8_io_out_activate),
    .io_out_weight(PE_Array_3_8_io_out_weight),
    .io_out_psum(PE_Array_3_8_io_out_psum)
  );
  basic_PE PE_Array_3_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_9_clock),
    .reset(PE_Array_3_9_reset),
    .io_in_activate(PE_Array_3_9_io_in_activate),
    .io_in_weight(PE_Array_3_9_io_in_weight),
    .io_in_psum(PE_Array_3_9_io_in_psum),
    .io_in_flow(PE_Array_3_9_io_in_flow),
    .io_in_shift(PE_Array_3_9_io_in_shift),
    .io_out_activate(PE_Array_3_9_io_out_activate),
    .io_out_weight(PE_Array_3_9_io_out_weight),
    .io_out_psum(PE_Array_3_9_io_out_psum)
  );
  basic_PE PE_Array_3_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_10_clock),
    .reset(PE_Array_3_10_reset),
    .io_in_activate(PE_Array_3_10_io_in_activate),
    .io_in_weight(PE_Array_3_10_io_in_weight),
    .io_in_psum(PE_Array_3_10_io_in_psum),
    .io_in_flow(PE_Array_3_10_io_in_flow),
    .io_in_shift(PE_Array_3_10_io_in_shift),
    .io_out_activate(PE_Array_3_10_io_out_activate),
    .io_out_weight(PE_Array_3_10_io_out_weight),
    .io_out_psum(PE_Array_3_10_io_out_psum)
  );
  basic_PE PE_Array_3_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_11_clock),
    .reset(PE_Array_3_11_reset),
    .io_in_activate(PE_Array_3_11_io_in_activate),
    .io_in_weight(PE_Array_3_11_io_in_weight),
    .io_in_psum(PE_Array_3_11_io_in_psum),
    .io_in_flow(PE_Array_3_11_io_in_flow),
    .io_in_shift(PE_Array_3_11_io_in_shift),
    .io_out_activate(PE_Array_3_11_io_out_activate),
    .io_out_weight(PE_Array_3_11_io_out_weight),
    .io_out_psum(PE_Array_3_11_io_out_psum)
  );
  basic_PE PE_Array_3_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_12_clock),
    .reset(PE_Array_3_12_reset),
    .io_in_activate(PE_Array_3_12_io_in_activate),
    .io_in_weight(PE_Array_3_12_io_in_weight),
    .io_in_psum(PE_Array_3_12_io_in_psum),
    .io_in_flow(PE_Array_3_12_io_in_flow),
    .io_in_shift(PE_Array_3_12_io_in_shift),
    .io_out_activate(PE_Array_3_12_io_out_activate),
    .io_out_weight(PE_Array_3_12_io_out_weight),
    .io_out_psum(PE_Array_3_12_io_out_psum)
  );
  basic_PE PE_Array_3_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_13_clock),
    .reset(PE_Array_3_13_reset),
    .io_in_activate(PE_Array_3_13_io_in_activate),
    .io_in_weight(PE_Array_3_13_io_in_weight),
    .io_in_psum(PE_Array_3_13_io_in_psum),
    .io_in_flow(PE_Array_3_13_io_in_flow),
    .io_in_shift(PE_Array_3_13_io_in_shift),
    .io_out_activate(PE_Array_3_13_io_out_activate),
    .io_out_weight(PE_Array_3_13_io_out_weight),
    .io_out_psum(PE_Array_3_13_io_out_psum)
  );
  basic_PE PE_Array_3_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_14_clock),
    .reset(PE_Array_3_14_reset),
    .io_in_activate(PE_Array_3_14_io_in_activate),
    .io_in_weight(PE_Array_3_14_io_in_weight),
    .io_in_psum(PE_Array_3_14_io_in_psum),
    .io_in_flow(PE_Array_3_14_io_in_flow),
    .io_in_shift(PE_Array_3_14_io_in_shift),
    .io_out_activate(PE_Array_3_14_io_out_activate),
    .io_out_weight(PE_Array_3_14_io_out_weight),
    .io_out_psum(PE_Array_3_14_io_out_psum)
  );
  basic_PE PE_Array_3_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_15_clock),
    .reset(PE_Array_3_15_reset),
    .io_in_activate(PE_Array_3_15_io_in_activate),
    .io_in_weight(PE_Array_3_15_io_in_weight),
    .io_in_psum(PE_Array_3_15_io_in_psum),
    .io_in_flow(PE_Array_3_15_io_in_flow),
    .io_in_shift(PE_Array_3_15_io_in_shift),
    .io_out_activate(PE_Array_3_15_io_out_activate),
    .io_out_weight(PE_Array_3_15_io_out_weight),
    .io_out_psum(PE_Array_3_15_io_out_psum)
  );
  basic_PE PE_Array_3_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_16_clock),
    .reset(PE_Array_3_16_reset),
    .io_in_activate(PE_Array_3_16_io_in_activate),
    .io_in_weight(PE_Array_3_16_io_in_weight),
    .io_in_psum(PE_Array_3_16_io_in_psum),
    .io_in_flow(PE_Array_3_16_io_in_flow),
    .io_in_shift(PE_Array_3_16_io_in_shift),
    .io_out_activate(PE_Array_3_16_io_out_activate),
    .io_out_weight(PE_Array_3_16_io_out_weight),
    .io_out_psum(PE_Array_3_16_io_out_psum)
  );
  basic_PE PE_Array_3_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_17_clock),
    .reset(PE_Array_3_17_reset),
    .io_in_activate(PE_Array_3_17_io_in_activate),
    .io_in_weight(PE_Array_3_17_io_in_weight),
    .io_in_psum(PE_Array_3_17_io_in_psum),
    .io_in_flow(PE_Array_3_17_io_in_flow),
    .io_in_shift(PE_Array_3_17_io_in_shift),
    .io_out_activate(PE_Array_3_17_io_out_activate),
    .io_out_weight(PE_Array_3_17_io_out_weight),
    .io_out_psum(PE_Array_3_17_io_out_psum)
  );
  basic_PE PE_Array_3_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_18_clock),
    .reset(PE_Array_3_18_reset),
    .io_in_activate(PE_Array_3_18_io_in_activate),
    .io_in_weight(PE_Array_3_18_io_in_weight),
    .io_in_psum(PE_Array_3_18_io_in_psum),
    .io_in_flow(PE_Array_3_18_io_in_flow),
    .io_in_shift(PE_Array_3_18_io_in_shift),
    .io_out_activate(PE_Array_3_18_io_out_activate),
    .io_out_weight(PE_Array_3_18_io_out_weight),
    .io_out_psum(PE_Array_3_18_io_out_psum)
  );
  basic_PE PE_Array_3_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_19_clock),
    .reset(PE_Array_3_19_reset),
    .io_in_activate(PE_Array_3_19_io_in_activate),
    .io_in_weight(PE_Array_3_19_io_in_weight),
    .io_in_psum(PE_Array_3_19_io_in_psum),
    .io_in_flow(PE_Array_3_19_io_in_flow),
    .io_in_shift(PE_Array_3_19_io_in_shift),
    .io_out_activate(PE_Array_3_19_io_out_activate),
    .io_out_weight(PE_Array_3_19_io_out_weight),
    .io_out_psum(PE_Array_3_19_io_out_psum)
  );
  basic_PE PE_Array_3_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_20_clock),
    .reset(PE_Array_3_20_reset),
    .io_in_activate(PE_Array_3_20_io_in_activate),
    .io_in_weight(PE_Array_3_20_io_in_weight),
    .io_in_psum(PE_Array_3_20_io_in_psum),
    .io_in_flow(PE_Array_3_20_io_in_flow),
    .io_in_shift(PE_Array_3_20_io_in_shift),
    .io_out_activate(PE_Array_3_20_io_out_activate),
    .io_out_weight(PE_Array_3_20_io_out_weight),
    .io_out_psum(PE_Array_3_20_io_out_psum)
  );
  basic_PE PE_Array_3_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_21_clock),
    .reset(PE_Array_3_21_reset),
    .io_in_activate(PE_Array_3_21_io_in_activate),
    .io_in_weight(PE_Array_3_21_io_in_weight),
    .io_in_psum(PE_Array_3_21_io_in_psum),
    .io_in_flow(PE_Array_3_21_io_in_flow),
    .io_in_shift(PE_Array_3_21_io_in_shift),
    .io_out_activate(PE_Array_3_21_io_out_activate),
    .io_out_weight(PE_Array_3_21_io_out_weight),
    .io_out_psum(PE_Array_3_21_io_out_psum)
  );
  basic_PE PE_Array_3_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_22_clock),
    .reset(PE_Array_3_22_reset),
    .io_in_activate(PE_Array_3_22_io_in_activate),
    .io_in_weight(PE_Array_3_22_io_in_weight),
    .io_in_psum(PE_Array_3_22_io_in_psum),
    .io_in_flow(PE_Array_3_22_io_in_flow),
    .io_in_shift(PE_Array_3_22_io_in_shift),
    .io_out_activate(PE_Array_3_22_io_out_activate),
    .io_out_weight(PE_Array_3_22_io_out_weight),
    .io_out_psum(PE_Array_3_22_io_out_psum)
  );
  basic_PE PE_Array_3_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_23_clock),
    .reset(PE_Array_3_23_reset),
    .io_in_activate(PE_Array_3_23_io_in_activate),
    .io_in_weight(PE_Array_3_23_io_in_weight),
    .io_in_psum(PE_Array_3_23_io_in_psum),
    .io_in_flow(PE_Array_3_23_io_in_flow),
    .io_in_shift(PE_Array_3_23_io_in_shift),
    .io_out_activate(PE_Array_3_23_io_out_activate),
    .io_out_weight(PE_Array_3_23_io_out_weight),
    .io_out_psum(PE_Array_3_23_io_out_psum)
  );
  basic_PE PE_Array_3_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_24_clock),
    .reset(PE_Array_3_24_reset),
    .io_in_activate(PE_Array_3_24_io_in_activate),
    .io_in_weight(PE_Array_3_24_io_in_weight),
    .io_in_psum(PE_Array_3_24_io_in_psum),
    .io_in_flow(PE_Array_3_24_io_in_flow),
    .io_in_shift(PE_Array_3_24_io_in_shift),
    .io_out_activate(PE_Array_3_24_io_out_activate),
    .io_out_weight(PE_Array_3_24_io_out_weight),
    .io_out_psum(PE_Array_3_24_io_out_psum)
  );
  basic_PE PE_Array_3_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_25_clock),
    .reset(PE_Array_3_25_reset),
    .io_in_activate(PE_Array_3_25_io_in_activate),
    .io_in_weight(PE_Array_3_25_io_in_weight),
    .io_in_psum(PE_Array_3_25_io_in_psum),
    .io_in_flow(PE_Array_3_25_io_in_flow),
    .io_in_shift(PE_Array_3_25_io_in_shift),
    .io_out_activate(PE_Array_3_25_io_out_activate),
    .io_out_weight(PE_Array_3_25_io_out_weight),
    .io_out_psum(PE_Array_3_25_io_out_psum)
  );
  basic_PE PE_Array_3_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_26_clock),
    .reset(PE_Array_3_26_reset),
    .io_in_activate(PE_Array_3_26_io_in_activate),
    .io_in_weight(PE_Array_3_26_io_in_weight),
    .io_in_psum(PE_Array_3_26_io_in_psum),
    .io_in_flow(PE_Array_3_26_io_in_flow),
    .io_in_shift(PE_Array_3_26_io_in_shift),
    .io_out_activate(PE_Array_3_26_io_out_activate),
    .io_out_weight(PE_Array_3_26_io_out_weight),
    .io_out_psum(PE_Array_3_26_io_out_psum)
  );
  basic_PE PE_Array_3_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_27_clock),
    .reset(PE_Array_3_27_reset),
    .io_in_activate(PE_Array_3_27_io_in_activate),
    .io_in_weight(PE_Array_3_27_io_in_weight),
    .io_in_psum(PE_Array_3_27_io_in_psum),
    .io_in_flow(PE_Array_3_27_io_in_flow),
    .io_in_shift(PE_Array_3_27_io_in_shift),
    .io_out_activate(PE_Array_3_27_io_out_activate),
    .io_out_weight(PE_Array_3_27_io_out_weight),
    .io_out_psum(PE_Array_3_27_io_out_psum)
  );
  basic_PE PE_Array_3_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_28_clock),
    .reset(PE_Array_3_28_reset),
    .io_in_activate(PE_Array_3_28_io_in_activate),
    .io_in_weight(PE_Array_3_28_io_in_weight),
    .io_in_psum(PE_Array_3_28_io_in_psum),
    .io_in_flow(PE_Array_3_28_io_in_flow),
    .io_in_shift(PE_Array_3_28_io_in_shift),
    .io_out_activate(PE_Array_3_28_io_out_activate),
    .io_out_weight(PE_Array_3_28_io_out_weight),
    .io_out_psum(PE_Array_3_28_io_out_psum)
  );
  basic_PE PE_Array_3_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_29_clock),
    .reset(PE_Array_3_29_reset),
    .io_in_activate(PE_Array_3_29_io_in_activate),
    .io_in_weight(PE_Array_3_29_io_in_weight),
    .io_in_psum(PE_Array_3_29_io_in_psum),
    .io_in_flow(PE_Array_3_29_io_in_flow),
    .io_in_shift(PE_Array_3_29_io_in_shift),
    .io_out_activate(PE_Array_3_29_io_out_activate),
    .io_out_weight(PE_Array_3_29_io_out_weight),
    .io_out_psum(PE_Array_3_29_io_out_psum)
  );
  basic_PE PE_Array_3_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_30_clock),
    .reset(PE_Array_3_30_reset),
    .io_in_activate(PE_Array_3_30_io_in_activate),
    .io_in_weight(PE_Array_3_30_io_in_weight),
    .io_in_psum(PE_Array_3_30_io_in_psum),
    .io_in_flow(PE_Array_3_30_io_in_flow),
    .io_in_shift(PE_Array_3_30_io_in_shift),
    .io_out_activate(PE_Array_3_30_io_out_activate),
    .io_out_weight(PE_Array_3_30_io_out_weight),
    .io_out_psum(PE_Array_3_30_io_out_psum)
  );
  basic_PE PE_Array_3_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_31_clock),
    .reset(PE_Array_3_31_reset),
    .io_in_activate(PE_Array_3_31_io_in_activate),
    .io_in_weight(PE_Array_3_31_io_in_weight),
    .io_in_psum(PE_Array_3_31_io_in_psum),
    .io_in_flow(PE_Array_3_31_io_in_flow),
    .io_in_shift(PE_Array_3_31_io_in_shift),
    .io_out_activate(PE_Array_3_31_io_out_activate),
    .io_out_weight(PE_Array_3_31_io_out_weight),
    .io_out_psum(PE_Array_3_31_io_out_psum)
  );
  basic_PE PE_Array_4_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_0_clock),
    .reset(PE_Array_4_0_reset),
    .io_in_activate(PE_Array_4_0_io_in_activate),
    .io_in_weight(PE_Array_4_0_io_in_weight),
    .io_in_psum(PE_Array_4_0_io_in_psum),
    .io_in_flow(PE_Array_4_0_io_in_flow),
    .io_in_shift(PE_Array_4_0_io_in_shift),
    .io_out_activate(PE_Array_4_0_io_out_activate),
    .io_out_weight(PE_Array_4_0_io_out_weight),
    .io_out_psum(PE_Array_4_0_io_out_psum)
  );
  basic_PE PE_Array_4_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_1_clock),
    .reset(PE_Array_4_1_reset),
    .io_in_activate(PE_Array_4_1_io_in_activate),
    .io_in_weight(PE_Array_4_1_io_in_weight),
    .io_in_psum(PE_Array_4_1_io_in_psum),
    .io_in_flow(PE_Array_4_1_io_in_flow),
    .io_in_shift(PE_Array_4_1_io_in_shift),
    .io_out_activate(PE_Array_4_1_io_out_activate),
    .io_out_weight(PE_Array_4_1_io_out_weight),
    .io_out_psum(PE_Array_4_1_io_out_psum)
  );
  basic_PE PE_Array_4_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_2_clock),
    .reset(PE_Array_4_2_reset),
    .io_in_activate(PE_Array_4_2_io_in_activate),
    .io_in_weight(PE_Array_4_2_io_in_weight),
    .io_in_psum(PE_Array_4_2_io_in_psum),
    .io_in_flow(PE_Array_4_2_io_in_flow),
    .io_in_shift(PE_Array_4_2_io_in_shift),
    .io_out_activate(PE_Array_4_2_io_out_activate),
    .io_out_weight(PE_Array_4_2_io_out_weight),
    .io_out_psum(PE_Array_4_2_io_out_psum)
  );
  basic_PE PE_Array_4_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_3_clock),
    .reset(PE_Array_4_3_reset),
    .io_in_activate(PE_Array_4_3_io_in_activate),
    .io_in_weight(PE_Array_4_3_io_in_weight),
    .io_in_psum(PE_Array_4_3_io_in_psum),
    .io_in_flow(PE_Array_4_3_io_in_flow),
    .io_in_shift(PE_Array_4_3_io_in_shift),
    .io_out_activate(PE_Array_4_3_io_out_activate),
    .io_out_weight(PE_Array_4_3_io_out_weight),
    .io_out_psum(PE_Array_4_3_io_out_psum)
  );
  basic_PE PE_Array_4_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_4_clock),
    .reset(PE_Array_4_4_reset),
    .io_in_activate(PE_Array_4_4_io_in_activate),
    .io_in_weight(PE_Array_4_4_io_in_weight),
    .io_in_psum(PE_Array_4_4_io_in_psum),
    .io_in_flow(PE_Array_4_4_io_in_flow),
    .io_in_shift(PE_Array_4_4_io_in_shift),
    .io_out_activate(PE_Array_4_4_io_out_activate),
    .io_out_weight(PE_Array_4_4_io_out_weight),
    .io_out_psum(PE_Array_4_4_io_out_psum)
  );
  basic_PE PE_Array_4_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_5_clock),
    .reset(PE_Array_4_5_reset),
    .io_in_activate(PE_Array_4_5_io_in_activate),
    .io_in_weight(PE_Array_4_5_io_in_weight),
    .io_in_psum(PE_Array_4_5_io_in_psum),
    .io_in_flow(PE_Array_4_5_io_in_flow),
    .io_in_shift(PE_Array_4_5_io_in_shift),
    .io_out_activate(PE_Array_4_5_io_out_activate),
    .io_out_weight(PE_Array_4_5_io_out_weight),
    .io_out_psum(PE_Array_4_5_io_out_psum)
  );
  basic_PE PE_Array_4_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_6_clock),
    .reset(PE_Array_4_6_reset),
    .io_in_activate(PE_Array_4_6_io_in_activate),
    .io_in_weight(PE_Array_4_6_io_in_weight),
    .io_in_psum(PE_Array_4_6_io_in_psum),
    .io_in_flow(PE_Array_4_6_io_in_flow),
    .io_in_shift(PE_Array_4_6_io_in_shift),
    .io_out_activate(PE_Array_4_6_io_out_activate),
    .io_out_weight(PE_Array_4_6_io_out_weight),
    .io_out_psum(PE_Array_4_6_io_out_psum)
  );
  basic_PE PE_Array_4_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_7_clock),
    .reset(PE_Array_4_7_reset),
    .io_in_activate(PE_Array_4_7_io_in_activate),
    .io_in_weight(PE_Array_4_7_io_in_weight),
    .io_in_psum(PE_Array_4_7_io_in_psum),
    .io_in_flow(PE_Array_4_7_io_in_flow),
    .io_in_shift(PE_Array_4_7_io_in_shift),
    .io_out_activate(PE_Array_4_7_io_out_activate),
    .io_out_weight(PE_Array_4_7_io_out_weight),
    .io_out_psum(PE_Array_4_7_io_out_psum)
  );
  basic_PE PE_Array_4_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_8_clock),
    .reset(PE_Array_4_8_reset),
    .io_in_activate(PE_Array_4_8_io_in_activate),
    .io_in_weight(PE_Array_4_8_io_in_weight),
    .io_in_psum(PE_Array_4_8_io_in_psum),
    .io_in_flow(PE_Array_4_8_io_in_flow),
    .io_in_shift(PE_Array_4_8_io_in_shift),
    .io_out_activate(PE_Array_4_8_io_out_activate),
    .io_out_weight(PE_Array_4_8_io_out_weight),
    .io_out_psum(PE_Array_4_8_io_out_psum)
  );
  basic_PE PE_Array_4_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_9_clock),
    .reset(PE_Array_4_9_reset),
    .io_in_activate(PE_Array_4_9_io_in_activate),
    .io_in_weight(PE_Array_4_9_io_in_weight),
    .io_in_psum(PE_Array_4_9_io_in_psum),
    .io_in_flow(PE_Array_4_9_io_in_flow),
    .io_in_shift(PE_Array_4_9_io_in_shift),
    .io_out_activate(PE_Array_4_9_io_out_activate),
    .io_out_weight(PE_Array_4_9_io_out_weight),
    .io_out_psum(PE_Array_4_9_io_out_psum)
  );
  basic_PE PE_Array_4_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_10_clock),
    .reset(PE_Array_4_10_reset),
    .io_in_activate(PE_Array_4_10_io_in_activate),
    .io_in_weight(PE_Array_4_10_io_in_weight),
    .io_in_psum(PE_Array_4_10_io_in_psum),
    .io_in_flow(PE_Array_4_10_io_in_flow),
    .io_in_shift(PE_Array_4_10_io_in_shift),
    .io_out_activate(PE_Array_4_10_io_out_activate),
    .io_out_weight(PE_Array_4_10_io_out_weight),
    .io_out_psum(PE_Array_4_10_io_out_psum)
  );
  basic_PE PE_Array_4_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_11_clock),
    .reset(PE_Array_4_11_reset),
    .io_in_activate(PE_Array_4_11_io_in_activate),
    .io_in_weight(PE_Array_4_11_io_in_weight),
    .io_in_psum(PE_Array_4_11_io_in_psum),
    .io_in_flow(PE_Array_4_11_io_in_flow),
    .io_in_shift(PE_Array_4_11_io_in_shift),
    .io_out_activate(PE_Array_4_11_io_out_activate),
    .io_out_weight(PE_Array_4_11_io_out_weight),
    .io_out_psum(PE_Array_4_11_io_out_psum)
  );
  basic_PE PE_Array_4_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_12_clock),
    .reset(PE_Array_4_12_reset),
    .io_in_activate(PE_Array_4_12_io_in_activate),
    .io_in_weight(PE_Array_4_12_io_in_weight),
    .io_in_psum(PE_Array_4_12_io_in_psum),
    .io_in_flow(PE_Array_4_12_io_in_flow),
    .io_in_shift(PE_Array_4_12_io_in_shift),
    .io_out_activate(PE_Array_4_12_io_out_activate),
    .io_out_weight(PE_Array_4_12_io_out_weight),
    .io_out_psum(PE_Array_4_12_io_out_psum)
  );
  basic_PE PE_Array_4_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_13_clock),
    .reset(PE_Array_4_13_reset),
    .io_in_activate(PE_Array_4_13_io_in_activate),
    .io_in_weight(PE_Array_4_13_io_in_weight),
    .io_in_psum(PE_Array_4_13_io_in_psum),
    .io_in_flow(PE_Array_4_13_io_in_flow),
    .io_in_shift(PE_Array_4_13_io_in_shift),
    .io_out_activate(PE_Array_4_13_io_out_activate),
    .io_out_weight(PE_Array_4_13_io_out_weight),
    .io_out_psum(PE_Array_4_13_io_out_psum)
  );
  basic_PE PE_Array_4_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_14_clock),
    .reset(PE_Array_4_14_reset),
    .io_in_activate(PE_Array_4_14_io_in_activate),
    .io_in_weight(PE_Array_4_14_io_in_weight),
    .io_in_psum(PE_Array_4_14_io_in_psum),
    .io_in_flow(PE_Array_4_14_io_in_flow),
    .io_in_shift(PE_Array_4_14_io_in_shift),
    .io_out_activate(PE_Array_4_14_io_out_activate),
    .io_out_weight(PE_Array_4_14_io_out_weight),
    .io_out_psum(PE_Array_4_14_io_out_psum)
  );
  basic_PE PE_Array_4_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_15_clock),
    .reset(PE_Array_4_15_reset),
    .io_in_activate(PE_Array_4_15_io_in_activate),
    .io_in_weight(PE_Array_4_15_io_in_weight),
    .io_in_psum(PE_Array_4_15_io_in_psum),
    .io_in_flow(PE_Array_4_15_io_in_flow),
    .io_in_shift(PE_Array_4_15_io_in_shift),
    .io_out_activate(PE_Array_4_15_io_out_activate),
    .io_out_weight(PE_Array_4_15_io_out_weight),
    .io_out_psum(PE_Array_4_15_io_out_psum)
  );
  basic_PE PE_Array_4_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_16_clock),
    .reset(PE_Array_4_16_reset),
    .io_in_activate(PE_Array_4_16_io_in_activate),
    .io_in_weight(PE_Array_4_16_io_in_weight),
    .io_in_psum(PE_Array_4_16_io_in_psum),
    .io_in_flow(PE_Array_4_16_io_in_flow),
    .io_in_shift(PE_Array_4_16_io_in_shift),
    .io_out_activate(PE_Array_4_16_io_out_activate),
    .io_out_weight(PE_Array_4_16_io_out_weight),
    .io_out_psum(PE_Array_4_16_io_out_psum)
  );
  basic_PE PE_Array_4_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_17_clock),
    .reset(PE_Array_4_17_reset),
    .io_in_activate(PE_Array_4_17_io_in_activate),
    .io_in_weight(PE_Array_4_17_io_in_weight),
    .io_in_psum(PE_Array_4_17_io_in_psum),
    .io_in_flow(PE_Array_4_17_io_in_flow),
    .io_in_shift(PE_Array_4_17_io_in_shift),
    .io_out_activate(PE_Array_4_17_io_out_activate),
    .io_out_weight(PE_Array_4_17_io_out_weight),
    .io_out_psum(PE_Array_4_17_io_out_psum)
  );
  basic_PE PE_Array_4_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_18_clock),
    .reset(PE_Array_4_18_reset),
    .io_in_activate(PE_Array_4_18_io_in_activate),
    .io_in_weight(PE_Array_4_18_io_in_weight),
    .io_in_psum(PE_Array_4_18_io_in_psum),
    .io_in_flow(PE_Array_4_18_io_in_flow),
    .io_in_shift(PE_Array_4_18_io_in_shift),
    .io_out_activate(PE_Array_4_18_io_out_activate),
    .io_out_weight(PE_Array_4_18_io_out_weight),
    .io_out_psum(PE_Array_4_18_io_out_psum)
  );
  basic_PE PE_Array_4_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_19_clock),
    .reset(PE_Array_4_19_reset),
    .io_in_activate(PE_Array_4_19_io_in_activate),
    .io_in_weight(PE_Array_4_19_io_in_weight),
    .io_in_psum(PE_Array_4_19_io_in_psum),
    .io_in_flow(PE_Array_4_19_io_in_flow),
    .io_in_shift(PE_Array_4_19_io_in_shift),
    .io_out_activate(PE_Array_4_19_io_out_activate),
    .io_out_weight(PE_Array_4_19_io_out_weight),
    .io_out_psum(PE_Array_4_19_io_out_psum)
  );
  basic_PE PE_Array_4_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_20_clock),
    .reset(PE_Array_4_20_reset),
    .io_in_activate(PE_Array_4_20_io_in_activate),
    .io_in_weight(PE_Array_4_20_io_in_weight),
    .io_in_psum(PE_Array_4_20_io_in_psum),
    .io_in_flow(PE_Array_4_20_io_in_flow),
    .io_in_shift(PE_Array_4_20_io_in_shift),
    .io_out_activate(PE_Array_4_20_io_out_activate),
    .io_out_weight(PE_Array_4_20_io_out_weight),
    .io_out_psum(PE_Array_4_20_io_out_psum)
  );
  basic_PE PE_Array_4_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_21_clock),
    .reset(PE_Array_4_21_reset),
    .io_in_activate(PE_Array_4_21_io_in_activate),
    .io_in_weight(PE_Array_4_21_io_in_weight),
    .io_in_psum(PE_Array_4_21_io_in_psum),
    .io_in_flow(PE_Array_4_21_io_in_flow),
    .io_in_shift(PE_Array_4_21_io_in_shift),
    .io_out_activate(PE_Array_4_21_io_out_activate),
    .io_out_weight(PE_Array_4_21_io_out_weight),
    .io_out_psum(PE_Array_4_21_io_out_psum)
  );
  basic_PE PE_Array_4_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_22_clock),
    .reset(PE_Array_4_22_reset),
    .io_in_activate(PE_Array_4_22_io_in_activate),
    .io_in_weight(PE_Array_4_22_io_in_weight),
    .io_in_psum(PE_Array_4_22_io_in_psum),
    .io_in_flow(PE_Array_4_22_io_in_flow),
    .io_in_shift(PE_Array_4_22_io_in_shift),
    .io_out_activate(PE_Array_4_22_io_out_activate),
    .io_out_weight(PE_Array_4_22_io_out_weight),
    .io_out_psum(PE_Array_4_22_io_out_psum)
  );
  basic_PE PE_Array_4_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_23_clock),
    .reset(PE_Array_4_23_reset),
    .io_in_activate(PE_Array_4_23_io_in_activate),
    .io_in_weight(PE_Array_4_23_io_in_weight),
    .io_in_psum(PE_Array_4_23_io_in_psum),
    .io_in_flow(PE_Array_4_23_io_in_flow),
    .io_in_shift(PE_Array_4_23_io_in_shift),
    .io_out_activate(PE_Array_4_23_io_out_activate),
    .io_out_weight(PE_Array_4_23_io_out_weight),
    .io_out_psum(PE_Array_4_23_io_out_psum)
  );
  basic_PE PE_Array_4_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_24_clock),
    .reset(PE_Array_4_24_reset),
    .io_in_activate(PE_Array_4_24_io_in_activate),
    .io_in_weight(PE_Array_4_24_io_in_weight),
    .io_in_psum(PE_Array_4_24_io_in_psum),
    .io_in_flow(PE_Array_4_24_io_in_flow),
    .io_in_shift(PE_Array_4_24_io_in_shift),
    .io_out_activate(PE_Array_4_24_io_out_activate),
    .io_out_weight(PE_Array_4_24_io_out_weight),
    .io_out_psum(PE_Array_4_24_io_out_psum)
  );
  basic_PE PE_Array_4_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_25_clock),
    .reset(PE_Array_4_25_reset),
    .io_in_activate(PE_Array_4_25_io_in_activate),
    .io_in_weight(PE_Array_4_25_io_in_weight),
    .io_in_psum(PE_Array_4_25_io_in_psum),
    .io_in_flow(PE_Array_4_25_io_in_flow),
    .io_in_shift(PE_Array_4_25_io_in_shift),
    .io_out_activate(PE_Array_4_25_io_out_activate),
    .io_out_weight(PE_Array_4_25_io_out_weight),
    .io_out_psum(PE_Array_4_25_io_out_psum)
  );
  basic_PE PE_Array_4_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_26_clock),
    .reset(PE_Array_4_26_reset),
    .io_in_activate(PE_Array_4_26_io_in_activate),
    .io_in_weight(PE_Array_4_26_io_in_weight),
    .io_in_psum(PE_Array_4_26_io_in_psum),
    .io_in_flow(PE_Array_4_26_io_in_flow),
    .io_in_shift(PE_Array_4_26_io_in_shift),
    .io_out_activate(PE_Array_4_26_io_out_activate),
    .io_out_weight(PE_Array_4_26_io_out_weight),
    .io_out_psum(PE_Array_4_26_io_out_psum)
  );
  basic_PE PE_Array_4_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_27_clock),
    .reset(PE_Array_4_27_reset),
    .io_in_activate(PE_Array_4_27_io_in_activate),
    .io_in_weight(PE_Array_4_27_io_in_weight),
    .io_in_psum(PE_Array_4_27_io_in_psum),
    .io_in_flow(PE_Array_4_27_io_in_flow),
    .io_in_shift(PE_Array_4_27_io_in_shift),
    .io_out_activate(PE_Array_4_27_io_out_activate),
    .io_out_weight(PE_Array_4_27_io_out_weight),
    .io_out_psum(PE_Array_4_27_io_out_psum)
  );
  basic_PE PE_Array_4_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_28_clock),
    .reset(PE_Array_4_28_reset),
    .io_in_activate(PE_Array_4_28_io_in_activate),
    .io_in_weight(PE_Array_4_28_io_in_weight),
    .io_in_psum(PE_Array_4_28_io_in_psum),
    .io_in_flow(PE_Array_4_28_io_in_flow),
    .io_in_shift(PE_Array_4_28_io_in_shift),
    .io_out_activate(PE_Array_4_28_io_out_activate),
    .io_out_weight(PE_Array_4_28_io_out_weight),
    .io_out_psum(PE_Array_4_28_io_out_psum)
  );
  basic_PE PE_Array_4_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_29_clock),
    .reset(PE_Array_4_29_reset),
    .io_in_activate(PE_Array_4_29_io_in_activate),
    .io_in_weight(PE_Array_4_29_io_in_weight),
    .io_in_psum(PE_Array_4_29_io_in_psum),
    .io_in_flow(PE_Array_4_29_io_in_flow),
    .io_in_shift(PE_Array_4_29_io_in_shift),
    .io_out_activate(PE_Array_4_29_io_out_activate),
    .io_out_weight(PE_Array_4_29_io_out_weight),
    .io_out_psum(PE_Array_4_29_io_out_psum)
  );
  basic_PE PE_Array_4_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_30_clock),
    .reset(PE_Array_4_30_reset),
    .io_in_activate(PE_Array_4_30_io_in_activate),
    .io_in_weight(PE_Array_4_30_io_in_weight),
    .io_in_psum(PE_Array_4_30_io_in_psum),
    .io_in_flow(PE_Array_4_30_io_in_flow),
    .io_in_shift(PE_Array_4_30_io_in_shift),
    .io_out_activate(PE_Array_4_30_io_out_activate),
    .io_out_weight(PE_Array_4_30_io_out_weight),
    .io_out_psum(PE_Array_4_30_io_out_psum)
  );
  basic_PE PE_Array_4_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_31_clock),
    .reset(PE_Array_4_31_reset),
    .io_in_activate(PE_Array_4_31_io_in_activate),
    .io_in_weight(PE_Array_4_31_io_in_weight),
    .io_in_psum(PE_Array_4_31_io_in_psum),
    .io_in_flow(PE_Array_4_31_io_in_flow),
    .io_in_shift(PE_Array_4_31_io_in_shift),
    .io_out_activate(PE_Array_4_31_io_out_activate),
    .io_out_weight(PE_Array_4_31_io_out_weight),
    .io_out_psum(PE_Array_4_31_io_out_psum)
  );
  basic_PE PE_Array_5_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_0_clock),
    .reset(PE_Array_5_0_reset),
    .io_in_activate(PE_Array_5_0_io_in_activate),
    .io_in_weight(PE_Array_5_0_io_in_weight),
    .io_in_psum(PE_Array_5_0_io_in_psum),
    .io_in_flow(PE_Array_5_0_io_in_flow),
    .io_in_shift(PE_Array_5_0_io_in_shift),
    .io_out_activate(PE_Array_5_0_io_out_activate),
    .io_out_weight(PE_Array_5_0_io_out_weight),
    .io_out_psum(PE_Array_5_0_io_out_psum)
  );
  basic_PE PE_Array_5_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_1_clock),
    .reset(PE_Array_5_1_reset),
    .io_in_activate(PE_Array_5_1_io_in_activate),
    .io_in_weight(PE_Array_5_1_io_in_weight),
    .io_in_psum(PE_Array_5_1_io_in_psum),
    .io_in_flow(PE_Array_5_1_io_in_flow),
    .io_in_shift(PE_Array_5_1_io_in_shift),
    .io_out_activate(PE_Array_5_1_io_out_activate),
    .io_out_weight(PE_Array_5_1_io_out_weight),
    .io_out_psum(PE_Array_5_1_io_out_psum)
  );
  basic_PE PE_Array_5_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_2_clock),
    .reset(PE_Array_5_2_reset),
    .io_in_activate(PE_Array_5_2_io_in_activate),
    .io_in_weight(PE_Array_5_2_io_in_weight),
    .io_in_psum(PE_Array_5_2_io_in_psum),
    .io_in_flow(PE_Array_5_2_io_in_flow),
    .io_in_shift(PE_Array_5_2_io_in_shift),
    .io_out_activate(PE_Array_5_2_io_out_activate),
    .io_out_weight(PE_Array_5_2_io_out_weight),
    .io_out_psum(PE_Array_5_2_io_out_psum)
  );
  basic_PE PE_Array_5_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_3_clock),
    .reset(PE_Array_5_3_reset),
    .io_in_activate(PE_Array_5_3_io_in_activate),
    .io_in_weight(PE_Array_5_3_io_in_weight),
    .io_in_psum(PE_Array_5_3_io_in_psum),
    .io_in_flow(PE_Array_5_3_io_in_flow),
    .io_in_shift(PE_Array_5_3_io_in_shift),
    .io_out_activate(PE_Array_5_3_io_out_activate),
    .io_out_weight(PE_Array_5_3_io_out_weight),
    .io_out_psum(PE_Array_5_3_io_out_psum)
  );
  basic_PE PE_Array_5_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_4_clock),
    .reset(PE_Array_5_4_reset),
    .io_in_activate(PE_Array_5_4_io_in_activate),
    .io_in_weight(PE_Array_5_4_io_in_weight),
    .io_in_psum(PE_Array_5_4_io_in_psum),
    .io_in_flow(PE_Array_5_4_io_in_flow),
    .io_in_shift(PE_Array_5_4_io_in_shift),
    .io_out_activate(PE_Array_5_4_io_out_activate),
    .io_out_weight(PE_Array_5_4_io_out_weight),
    .io_out_psum(PE_Array_5_4_io_out_psum)
  );
  basic_PE PE_Array_5_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_5_clock),
    .reset(PE_Array_5_5_reset),
    .io_in_activate(PE_Array_5_5_io_in_activate),
    .io_in_weight(PE_Array_5_5_io_in_weight),
    .io_in_psum(PE_Array_5_5_io_in_psum),
    .io_in_flow(PE_Array_5_5_io_in_flow),
    .io_in_shift(PE_Array_5_5_io_in_shift),
    .io_out_activate(PE_Array_5_5_io_out_activate),
    .io_out_weight(PE_Array_5_5_io_out_weight),
    .io_out_psum(PE_Array_5_5_io_out_psum)
  );
  basic_PE PE_Array_5_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_6_clock),
    .reset(PE_Array_5_6_reset),
    .io_in_activate(PE_Array_5_6_io_in_activate),
    .io_in_weight(PE_Array_5_6_io_in_weight),
    .io_in_psum(PE_Array_5_6_io_in_psum),
    .io_in_flow(PE_Array_5_6_io_in_flow),
    .io_in_shift(PE_Array_5_6_io_in_shift),
    .io_out_activate(PE_Array_5_6_io_out_activate),
    .io_out_weight(PE_Array_5_6_io_out_weight),
    .io_out_psum(PE_Array_5_6_io_out_psum)
  );
  basic_PE PE_Array_5_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_7_clock),
    .reset(PE_Array_5_7_reset),
    .io_in_activate(PE_Array_5_7_io_in_activate),
    .io_in_weight(PE_Array_5_7_io_in_weight),
    .io_in_psum(PE_Array_5_7_io_in_psum),
    .io_in_flow(PE_Array_5_7_io_in_flow),
    .io_in_shift(PE_Array_5_7_io_in_shift),
    .io_out_activate(PE_Array_5_7_io_out_activate),
    .io_out_weight(PE_Array_5_7_io_out_weight),
    .io_out_psum(PE_Array_5_7_io_out_psum)
  );
  basic_PE PE_Array_5_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_8_clock),
    .reset(PE_Array_5_8_reset),
    .io_in_activate(PE_Array_5_8_io_in_activate),
    .io_in_weight(PE_Array_5_8_io_in_weight),
    .io_in_psum(PE_Array_5_8_io_in_psum),
    .io_in_flow(PE_Array_5_8_io_in_flow),
    .io_in_shift(PE_Array_5_8_io_in_shift),
    .io_out_activate(PE_Array_5_8_io_out_activate),
    .io_out_weight(PE_Array_5_8_io_out_weight),
    .io_out_psum(PE_Array_5_8_io_out_psum)
  );
  basic_PE PE_Array_5_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_9_clock),
    .reset(PE_Array_5_9_reset),
    .io_in_activate(PE_Array_5_9_io_in_activate),
    .io_in_weight(PE_Array_5_9_io_in_weight),
    .io_in_psum(PE_Array_5_9_io_in_psum),
    .io_in_flow(PE_Array_5_9_io_in_flow),
    .io_in_shift(PE_Array_5_9_io_in_shift),
    .io_out_activate(PE_Array_5_9_io_out_activate),
    .io_out_weight(PE_Array_5_9_io_out_weight),
    .io_out_psum(PE_Array_5_9_io_out_psum)
  );
  basic_PE PE_Array_5_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_10_clock),
    .reset(PE_Array_5_10_reset),
    .io_in_activate(PE_Array_5_10_io_in_activate),
    .io_in_weight(PE_Array_5_10_io_in_weight),
    .io_in_psum(PE_Array_5_10_io_in_psum),
    .io_in_flow(PE_Array_5_10_io_in_flow),
    .io_in_shift(PE_Array_5_10_io_in_shift),
    .io_out_activate(PE_Array_5_10_io_out_activate),
    .io_out_weight(PE_Array_5_10_io_out_weight),
    .io_out_psum(PE_Array_5_10_io_out_psum)
  );
  basic_PE PE_Array_5_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_11_clock),
    .reset(PE_Array_5_11_reset),
    .io_in_activate(PE_Array_5_11_io_in_activate),
    .io_in_weight(PE_Array_5_11_io_in_weight),
    .io_in_psum(PE_Array_5_11_io_in_psum),
    .io_in_flow(PE_Array_5_11_io_in_flow),
    .io_in_shift(PE_Array_5_11_io_in_shift),
    .io_out_activate(PE_Array_5_11_io_out_activate),
    .io_out_weight(PE_Array_5_11_io_out_weight),
    .io_out_psum(PE_Array_5_11_io_out_psum)
  );
  basic_PE PE_Array_5_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_12_clock),
    .reset(PE_Array_5_12_reset),
    .io_in_activate(PE_Array_5_12_io_in_activate),
    .io_in_weight(PE_Array_5_12_io_in_weight),
    .io_in_psum(PE_Array_5_12_io_in_psum),
    .io_in_flow(PE_Array_5_12_io_in_flow),
    .io_in_shift(PE_Array_5_12_io_in_shift),
    .io_out_activate(PE_Array_5_12_io_out_activate),
    .io_out_weight(PE_Array_5_12_io_out_weight),
    .io_out_psum(PE_Array_5_12_io_out_psum)
  );
  basic_PE PE_Array_5_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_13_clock),
    .reset(PE_Array_5_13_reset),
    .io_in_activate(PE_Array_5_13_io_in_activate),
    .io_in_weight(PE_Array_5_13_io_in_weight),
    .io_in_psum(PE_Array_5_13_io_in_psum),
    .io_in_flow(PE_Array_5_13_io_in_flow),
    .io_in_shift(PE_Array_5_13_io_in_shift),
    .io_out_activate(PE_Array_5_13_io_out_activate),
    .io_out_weight(PE_Array_5_13_io_out_weight),
    .io_out_psum(PE_Array_5_13_io_out_psum)
  );
  basic_PE PE_Array_5_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_14_clock),
    .reset(PE_Array_5_14_reset),
    .io_in_activate(PE_Array_5_14_io_in_activate),
    .io_in_weight(PE_Array_5_14_io_in_weight),
    .io_in_psum(PE_Array_5_14_io_in_psum),
    .io_in_flow(PE_Array_5_14_io_in_flow),
    .io_in_shift(PE_Array_5_14_io_in_shift),
    .io_out_activate(PE_Array_5_14_io_out_activate),
    .io_out_weight(PE_Array_5_14_io_out_weight),
    .io_out_psum(PE_Array_5_14_io_out_psum)
  );
  basic_PE PE_Array_5_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_15_clock),
    .reset(PE_Array_5_15_reset),
    .io_in_activate(PE_Array_5_15_io_in_activate),
    .io_in_weight(PE_Array_5_15_io_in_weight),
    .io_in_psum(PE_Array_5_15_io_in_psum),
    .io_in_flow(PE_Array_5_15_io_in_flow),
    .io_in_shift(PE_Array_5_15_io_in_shift),
    .io_out_activate(PE_Array_5_15_io_out_activate),
    .io_out_weight(PE_Array_5_15_io_out_weight),
    .io_out_psum(PE_Array_5_15_io_out_psum)
  );
  basic_PE PE_Array_5_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_16_clock),
    .reset(PE_Array_5_16_reset),
    .io_in_activate(PE_Array_5_16_io_in_activate),
    .io_in_weight(PE_Array_5_16_io_in_weight),
    .io_in_psum(PE_Array_5_16_io_in_psum),
    .io_in_flow(PE_Array_5_16_io_in_flow),
    .io_in_shift(PE_Array_5_16_io_in_shift),
    .io_out_activate(PE_Array_5_16_io_out_activate),
    .io_out_weight(PE_Array_5_16_io_out_weight),
    .io_out_psum(PE_Array_5_16_io_out_psum)
  );
  basic_PE PE_Array_5_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_17_clock),
    .reset(PE_Array_5_17_reset),
    .io_in_activate(PE_Array_5_17_io_in_activate),
    .io_in_weight(PE_Array_5_17_io_in_weight),
    .io_in_psum(PE_Array_5_17_io_in_psum),
    .io_in_flow(PE_Array_5_17_io_in_flow),
    .io_in_shift(PE_Array_5_17_io_in_shift),
    .io_out_activate(PE_Array_5_17_io_out_activate),
    .io_out_weight(PE_Array_5_17_io_out_weight),
    .io_out_psum(PE_Array_5_17_io_out_psum)
  );
  basic_PE PE_Array_5_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_18_clock),
    .reset(PE_Array_5_18_reset),
    .io_in_activate(PE_Array_5_18_io_in_activate),
    .io_in_weight(PE_Array_5_18_io_in_weight),
    .io_in_psum(PE_Array_5_18_io_in_psum),
    .io_in_flow(PE_Array_5_18_io_in_flow),
    .io_in_shift(PE_Array_5_18_io_in_shift),
    .io_out_activate(PE_Array_5_18_io_out_activate),
    .io_out_weight(PE_Array_5_18_io_out_weight),
    .io_out_psum(PE_Array_5_18_io_out_psum)
  );
  basic_PE PE_Array_5_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_19_clock),
    .reset(PE_Array_5_19_reset),
    .io_in_activate(PE_Array_5_19_io_in_activate),
    .io_in_weight(PE_Array_5_19_io_in_weight),
    .io_in_psum(PE_Array_5_19_io_in_psum),
    .io_in_flow(PE_Array_5_19_io_in_flow),
    .io_in_shift(PE_Array_5_19_io_in_shift),
    .io_out_activate(PE_Array_5_19_io_out_activate),
    .io_out_weight(PE_Array_5_19_io_out_weight),
    .io_out_psum(PE_Array_5_19_io_out_psum)
  );
  basic_PE PE_Array_5_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_20_clock),
    .reset(PE_Array_5_20_reset),
    .io_in_activate(PE_Array_5_20_io_in_activate),
    .io_in_weight(PE_Array_5_20_io_in_weight),
    .io_in_psum(PE_Array_5_20_io_in_psum),
    .io_in_flow(PE_Array_5_20_io_in_flow),
    .io_in_shift(PE_Array_5_20_io_in_shift),
    .io_out_activate(PE_Array_5_20_io_out_activate),
    .io_out_weight(PE_Array_5_20_io_out_weight),
    .io_out_psum(PE_Array_5_20_io_out_psum)
  );
  basic_PE PE_Array_5_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_21_clock),
    .reset(PE_Array_5_21_reset),
    .io_in_activate(PE_Array_5_21_io_in_activate),
    .io_in_weight(PE_Array_5_21_io_in_weight),
    .io_in_psum(PE_Array_5_21_io_in_psum),
    .io_in_flow(PE_Array_5_21_io_in_flow),
    .io_in_shift(PE_Array_5_21_io_in_shift),
    .io_out_activate(PE_Array_5_21_io_out_activate),
    .io_out_weight(PE_Array_5_21_io_out_weight),
    .io_out_psum(PE_Array_5_21_io_out_psum)
  );
  basic_PE PE_Array_5_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_22_clock),
    .reset(PE_Array_5_22_reset),
    .io_in_activate(PE_Array_5_22_io_in_activate),
    .io_in_weight(PE_Array_5_22_io_in_weight),
    .io_in_psum(PE_Array_5_22_io_in_psum),
    .io_in_flow(PE_Array_5_22_io_in_flow),
    .io_in_shift(PE_Array_5_22_io_in_shift),
    .io_out_activate(PE_Array_5_22_io_out_activate),
    .io_out_weight(PE_Array_5_22_io_out_weight),
    .io_out_psum(PE_Array_5_22_io_out_psum)
  );
  basic_PE PE_Array_5_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_23_clock),
    .reset(PE_Array_5_23_reset),
    .io_in_activate(PE_Array_5_23_io_in_activate),
    .io_in_weight(PE_Array_5_23_io_in_weight),
    .io_in_psum(PE_Array_5_23_io_in_psum),
    .io_in_flow(PE_Array_5_23_io_in_flow),
    .io_in_shift(PE_Array_5_23_io_in_shift),
    .io_out_activate(PE_Array_5_23_io_out_activate),
    .io_out_weight(PE_Array_5_23_io_out_weight),
    .io_out_psum(PE_Array_5_23_io_out_psum)
  );
  basic_PE PE_Array_5_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_24_clock),
    .reset(PE_Array_5_24_reset),
    .io_in_activate(PE_Array_5_24_io_in_activate),
    .io_in_weight(PE_Array_5_24_io_in_weight),
    .io_in_psum(PE_Array_5_24_io_in_psum),
    .io_in_flow(PE_Array_5_24_io_in_flow),
    .io_in_shift(PE_Array_5_24_io_in_shift),
    .io_out_activate(PE_Array_5_24_io_out_activate),
    .io_out_weight(PE_Array_5_24_io_out_weight),
    .io_out_psum(PE_Array_5_24_io_out_psum)
  );
  basic_PE PE_Array_5_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_25_clock),
    .reset(PE_Array_5_25_reset),
    .io_in_activate(PE_Array_5_25_io_in_activate),
    .io_in_weight(PE_Array_5_25_io_in_weight),
    .io_in_psum(PE_Array_5_25_io_in_psum),
    .io_in_flow(PE_Array_5_25_io_in_flow),
    .io_in_shift(PE_Array_5_25_io_in_shift),
    .io_out_activate(PE_Array_5_25_io_out_activate),
    .io_out_weight(PE_Array_5_25_io_out_weight),
    .io_out_psum(PE_Array_5_25_io_out_psum)
  );
  basic_PE PE_Array_5_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_26_clock),
    .reset(PE_Array_5_26_reset),
    .io_in_activate(PE_Array_5_26_io_in_activate),
    .io_in_weight(PE_Array_5_26_io_in_weight),
    .io_in_psum(PE_Array_5_26_io_in_psum),
    .io_in_flow(PE_Array_5_26_io_in_flow),
    .io_in_shift(PE_Array_5_26_io_in_shift),
    .io_out_activate(PE_Array_5_26_io_out_activate),
    .io_out_weight(PE_Array_5_26_io_out_weight),
    .io_out_psum(PE_Array_5_26_io_out_psum)
  );
  basic_PE PE_Array_5_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_27_clock),
    .reset(PE_Array_5_27_reset),
    .io_in_activate(PE_Array_5_27_io_in_activate),
    .io_in_weight(PE_Array_5_27_io_in_weight),
    .io_in_psum(PE_Array_5_27_io_in_psum),
    .io_in_flow(PE_Array_5_27_io_in_flow),
    .io_in_shift(PE_Array_5_27_io_in_shift),
    .io_out_activate(PE_Array_5_27_io_out_activate),
    .io_out_weight(PE_Array_5_27_io_out_weight),
    .io_out_psum(PE_Array_5_27_io_out_psum)
  );
  basic_PE PE_Array_5_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_28_clock),
    .reset(PE_Array_5_28_reset),
    .io_in_activate(PE_Array_5_28_io_in_activate),
    .io_in_weight(PE_Array_5_28_io_in_weight),
    .io_in_psum(PE_Array_5_28_io_in_psum),
    .io_in_flow(PE_Array_5_28_io_in_flow),
    .io_in_shift(PE_Array_5_28_io_in_shift),
    .io_out_activate(PE_Array_5_28_io_out_activate),
    .io_out_weight(PE_Array_5_28_io_out_weight),
    .io_out_psum(PE_Array_5_28_io_out_psum)
  );
  basic_PE PE_Array_5_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_29_clock),
    .reset(PE_Array_5_29_reset),
    .io_in_activate(PE_Array_5_29_io_in_activate),
    .io_in_weight(PE_Array_5_29_io_in_weight),
    .io_in_psum(PE_Array_5_29_io_in_psum),
    .io_in_flow(PE_Array_5_29_io_in_flow),
    .io_in_shift(PE_Array_5_29_io_in_shift),
    .io_out_activate(PE_Array_5_29_io_out_activate),
    .io_out_weight(PE_Array_5_29_io_out_weight),
    .io_out_psum(PE_Array_5_29_io_out_psum)
  );
  basic_PE PE_Array_5_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_30_clock),
    .reset(PE_Array_5_30_reset),
    .io_in_activate(PE_Array_5_30_io_in_activate),
    .io_in_weight(PE_Array_5_30_io_in_weight),
    .io_in_psum(PE_Array_5_30_io_in_psum),
    .io_in_flow(PE_Array_5_30_io_in_flow),
    .io_in_shift(PE_Array_5_30_io_in_shift),
    .io_out_activate(PE_Array_5_30_io_out_activate),
    .io_out_weight(PE_Array_5_30_io_out_weight),
    .io_out_psum(PE_Array_5_30_io_out_psum)
  );
  basic_PE PE_Array_5_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_31_clock),
    .reset(PE_Array_5_31_reset),
    .io_in_activate(PE_Array_5_31_io_in_activate),
    .io_in_weight(PE_Array_5_31_io_in_weight),
    .io_in_psum(PE_Array_5_31_io_in_psum),
    .io_in_flow(PE_Array_5_31_io_in_flow),
    .io_in_shift(PE_Array_5_31_io_in_shift),
    .io_out_activate(PE_Array_5_31_io_out_activate),
    .io_out_weight(PE_Array_5_31_io_out_weight),
    .io_out_psum(PE_Array_5_31_io_out_psum)
  );
  basic_PE PE_Array_6_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_0_clock),
    .reset(PE_Array_6_0_reset),
    .io_in_activate(PE_Array_6_0_io_in_activate),
    .io_in_weight(PE_Array_6_0_io_in_weight),
    .io_in_psum(PE_Array_6_0_io_in_psum),
    .io_in_flow(PE_Array_6_0_io_in_flow),
    .io_in_shift(PE_Array_6_0_io_in_shift),
    .io_out_activate(PE_Array_6_0_io_out_activate),
    .io_out_weight(PE_Array_6_0_io_out_weight),
    .io_out_psum(PE_Array_6_0_io_out_psum)
  );
  basic_PE PE_Array_6_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_1_clock),
    .reset(PE_Array_6_1_reset),
    .io_in_activate(PE_Array_6_1_io_in_activate),
    .io_in_weight(PE_Array_6_1_io_in_weight),
    .io_in_psum(PE_Array_6_1_io_in_psum),
    .io_in_flow(PE_Array_6_1_io_in_flow),
    .io_in_shift(PE_Array_6_1_io_in_shift),
    .io_out_activate(PE_Array_6_1_io_out_activate),
    .io_out_weight(PE_Array_6_1_io_out_weight),
    .io_out_psum(PE_Array_6_1_io_out_psum)
  );
  basic_PE PE_Array_6_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_2_clock),
    .reset(PE_Array_6_2_reset),
    .io_in_activate(PE_Array_6_2_io_in_activate),
    .io_in_weight(PE_Array_6_2_io_in_weight),
    .io_in_psum(PE_Array_6_2_io_in_psum),
    .io_in_flow(PE_Array_6_2_io_in_flow),
    .io_in_shift(PE_Array_6_2_io_in_shift),
    .io_out_activate(PE_Array_6_2_io_out_activate),
    .io_out_weight(PE_Array_6_2_io_out_weight),
    .io_out_psum(PE_Array_6_2_io_out_psum)
  );
  basic_PE PE_Array_6_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_3_clock),
    .reset(PE_Array_6_3_reset),
    .io_in_activate(PE_Array_6_3_io_in_activate),
    .io_in_weight(PE_Array_6_3_io_in_weight),
    .io_in_psum(PE_Array_6_3_io_in_psum),
    .io_in_flow(PE_Array_6_3_io_in_flow),
    .io_in_shift(PE_Array_6_3_io_in_shift),
    .io_out_activate(PE_Array_6_3_io_out_activate),
    .io_out_weight(PE_Array_6_3_io_out_weight),
    .io_out_psum(PE_Array_6_3_io_out_psum)
  );
  basic_PE PE_Array_6_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_4_clock),
    .reset(PE_Array_6_4_reset),
    .io_in_activate(PE_Array_6_4_io_in_activate),
    .io_in_weight(PE_Array_6_4_io_in_weight),
    .io_in_psum(PE_Array_6_4_io_in_psum),
    .io_in_flow(PE_Array_6_4_io_in_flow),
    .io_in_shift(PE_Array_6_4_io_in_shift),
    .io_out_activate(PE_Array_6_4_io_out_activate),
    .io_out_weight(PE_Array_6_4_io_out_weight),
    .io_out_psum(PE_Array_6_4_io_out_psum)
  );
  basic_PE PE_Array_6_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_5_clock),
    .reset(PE_Array_6_5_reset),
    .io_in_activate(PE_Array_6_5_io_in_activate),
    .io_in_weight(PE_Array_6_5_io_in_weight),
    .io_in_psum(PE_Array_6_5_io_in_psum),
    .io_in_flow(PE_Array_6_5_io_in_flow),
    .io_in_shift(PE_Array_6_5_io_in_shift),
    .io_out_activate(PE_Array_6_5_io_out_activate),
    .io_out_weight(PE_Array_6_5_io_out_weight),
    .io_out_psum(PE_Array_6_5_io_out_psum)
  );
  basic_PE PE_Array_6_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_6_clock),
    .reset(PE_Array_6_6_reset),
    .io_in_activate(PE_Array_6_6_io_in_activate),
    .io_in_weight(PE_Array_6_6_io_in_weight),
    .io_in_psum(PE_Array_6_6_io_in_psum),
    .io_in_flow(PE_Array_6_6_io_in_flow),
    .io_in_shift(PE_Array_6_6_io_in_shift),
    .io_out_activate(PE_Array_6_6_io_out_activate),
    .io_out_weight(PE_Array_6_6_io_out_weight),
    .io_out_psum(PE_Array_6_6_io_out_psum)
  );
  basic_PE PE_Array_6_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_7_clock),
    .reset(PE_Array_6_7_reset),
    .io_in_activate(PE_Array_6_7_io_in_activate),
    .io_in_weight(PE_Array_6_7_io_in_weight),
    .io_in_psum(PE_Array_6_7_io_in_psum),
    .io_in_flow(PE_Array_6_7_io_in_flow),
    .io_in_shift(PE_Array_6_7_io_in_shift),
    .io_out_activate(PE_Array_6_7_io_out_activate),
    .io_out_weight(PE_Array_6_7_io_out_weight),
    .io_out_psum(PE_Array_6_7_io_out_psum)
  );
  basic_PE PE_Array_6_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_8_clock),
    .reset(PE_Array_6_8_reset),
    .io_in_activate(PE_Array_6_8_io_in_activate),
    .io_in_weight(PE_Array_6_8_io_in_weight),
    .io_in_psum(PE_Array_6_8_io_in_psum),
    .io_in_flow(PE_Array_6_8_io_in_flow),
    .io_in_shift(PE_Array_6_8_io_in_shift),
    .io_out_activate(PE_Array_6_8_io_out_activate),
    .io_out_weight(PE_Array_6_8_io_out_weight),
    .io_out_psum(PE_Array_6_8_io_out_psum)
  );
  basic_PE PE_Array_6_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_9_clock),
    .reset(PE_Array_6_9_reset),
    .io_in_activate(PE_Array_6_9_io_in_activate),
    .io_in_weight(PE_Array_6_9_io_in_weight),
    .io_in_psum(PE_Array_6_9_io_in_psum),
    .io_in_flow(PE_Array_6_9_io_in_flow),
    .io_in_shift(PE_Array_6_9_io_in_shift),
    .io_out_activate(PE_Array_6_9_io_out_activate),
    .io_out_weight(PE_Array_6_9_io_out_weight),
    .io_out_psum(PE_Array_6_9_io_out_psum)
  );
  basic_PE PE_Array_6_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_10_clock),
    .reset(PE_Array_6_10_reset),
    .io_in_activate(PE_Array_6_10_io_in_activate),
    .io_in_weight(PE_Array_6_10_io_in_weight),
    .io_in_psum(PE_Array_6_10_io_in_psum),
    .io_in_flow(PE_Array_6_10_io_in_flow),
    .io_in_shift(PE_Array_6_10_io_in_shift),
    .io_out_activate(PE_Array_6_10_io_out_activate),
    .io_out_weight(PE_Array_6_10_io_out_weight),
    .io_out_psum(PE_Array_6_10_io_out_psum)
  );
  basic_PE PE_Array_6_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_11_clock),
    .reset(PE_Array_6_11_reset),
    .io_in_activate(PE_Array_6_11_io_in_activate),
    .io_in_weight(PE_Array_6_11_io_in_weight),
    .io_in_psum(PE_Array_6_11_io_in_psum),
    .io_in_flow(PE_Array_6_11_io_in_flow),
    .io_in_shift(PE_Array_6_11_io_in_shift),
    .io_out_activate(PE_Array_6_11_io_out_activate),
    .io_out_weight(PE_Array_6_11_io_out_weight),
    .io_out_psum(PE_Array_6_11_io_out_psum)
  );
  basic_PE PE_Array_6_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_12_clock),
    .reset(PE_Array_6_12_reset),
    .io_in_activate(PE_Array_6_12_io_in_activate),
    .io_in_weight(PE_Array_6_12_io_in_weight),
    .io_in_psum(PE_Array_6_12_io_in_psum),
    .io_in_flow(PE_Array_6_12_io_in_flow),
    .io_in_shift(PE_Array_6_12_io_in_shift),
    .io_out_activate(PE_Array_6_12_io_out_activate),
    .io_out_weight(PE_Array_6_12_io_out_weight),
    .io_out_psum(PE_Array_6_12_io_out_psum)
  );
  basic_PE PE_Array_6_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_13_clock),
    .reset(PE_Array_6_13_reset),
    .io_in_activate(PE_Array_6_13_io_in_activate),
    .io_in_weight(PE_Array_6_13_io_in_weight),
    .io_in_psum(PE_Array_6_13_io_in_psum),
    .io_in_flow(PE_Array_6_13_io_in_flow),
    .io_in_shift(PE_Array_6_13_io_in_shift),
    .io_out_activate(PE_Array_6_13_io_out_activate),
    .io_out_weight(PE_Array_6_13_io_out_weight),
    .io_out_psum(PE_Array_6_13_io_out_psum)
  );
  basic_PE PE_Array_6_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_14_clock),
    .reset(PE_Array_6_14_reset),
    .io_in_activate(PE_Array_6_14_io_in_activate),
    .io_in_weight(PE_Array_6_14_io_in_weight),
    .io_in_psum(PE_Array_6_14_io_in_psum),
    .io_in_flow(PE_Array_6_14_io_in_flow),
    .io_in_shift(PE_Array_6_14_io_in_shift),
    .io_out_activate(PE_Array_6_14_io_out_activate),
    .io_out_weight(PE_Array_6_14_io_out_weight),
    .io_out_psum(PE_Array_6_14_io_out_psum)
  );
  basic_PE PE_Array_6_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_15_clock),
    .reset(PE_Array_6_15_reset),
    .io_in_activate(PE_Array_6_15_io_in_activate),
    .io_in_weight(PE_Array_6_15_io_in_weight),
    .io_in_psum(PE_Array_6_15_io_in_psum),
    .io_in_flow(PE_Array_6_15_io_in_flow),
    .io_in_shift(PE_Array_6_15_io_in_shift),
    .io_out_activate(PE_Array_6_15_io_out_activate),
    .io_out_weight(PE_Array_6_15_io_out_weight),
    .io_out_psum(PE_Array_6_15_io_out_psum)
  );
  basic_PE PE_Array_6_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_16_clock),
    .reset(PE_Array_6_16_reset),
    .io_in_activate(PE_Array_6_16_io_in_activate),
    .io_in_weight(PE_Array_6_16_io_in_weight),
    .io_in_psum(PE_Array_6_16_io_in_psum),
    .io_in_flow(PE_Array_6_16_io_in_flow),
    .io_in_shift(PE_Array_6_16_io_in_shift),
    .io_out_activate(PE_Array_6_16_io_out_activate),
    .io_out_weight(PE_Array_6_16_io_out_weight),
    .io_out_psum(PE_Array_6_16_io_out_psum)
  );
  basic_PE PE_Array_6_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_17_clock),
    .reset(PE_Array_6_17_reset),
    .io_in_activate(PE_Array_6_17_io_in_activate),
    .io_in_weight(PE_Array_6_17_io_in_weight),
    .io_in_psum(PE_Array_6_17_io_in_psum),
    .io_in_flow(PE_Array_6_17_io_in_flow),
    .io_in_shift(PE_Array_6_17_io_in_shift),
    .io_out_activate(PE_Array_6_17_io_out_activate),
    .io_out_weight(PE_Array_6_17_io_out_weight),
    .io_out_psum(PE_Array_6_17_io_out_psum)
  );
  basic_PE PE_Array_6_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_18_clock),
    .reset(PE_Array_6_18_reset),
    .io_in_activate(PE_Array_6_18_io_in_activate),
    .io_in_weight(PE_Array_6_18_io_in_weight),
    .io_in_psum(PE_Array_6_18_io_in_psum),
    .io_in_flow(PE_Array_6_18_io_in_flow),
    .io_in_shift(PE_Array_6_18_io_in_shift),
    .io_out_activate(PE_Array_6_18_io_out_activate),
    .io_out_weight(PE_Array_6_18_io_out_weight),
    .io_out_psum(PE_Array_6_18_io_out_psum)
  );
  basic_PE PE_Array_6_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_19_clock),
    .reset(PE_Array_6_19_reset),
    .io_in_activate(PE_Array_6_19_io_in_activate),
    .io_in_weight(PE_Array_6_19_io_in_weight),
    .io_in_psum(PE_Array_6_19_io_in_psum),
    .io_in_flow(PE_Array_6_19_io_in_flow),
    .io_in_shift(PE_Array_6_19_io_in_shift),
    .io_out_activate(PE_Array_6_19_io_out_activate),
    .io_out_weight(PE_Array_6_19_io_out_weight),
    .io_out_psum(PE_Array_6_19_io_out_psum)
  );
  basic_PE PE_Array_6_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_20_clock),
    .reset(PE_Array_6_20_reset),
    .io_in_activate(PE_Array_6_20_io_in_activate),
    .io_in_weight(PE_Array_6_20_io_in_weight),
    .io_in_psum(PE_Array_6_20_io_in_psum),
    .io_in_flow(PE_Array_6_20_io_in_flow),
    .io_in_shift(PE_Array_6_20_io_in_shift),
    .io_out_activate(PE_Array_6_20_io_out_activate),
    .io_out_weight(PE_Array_6_20_io_out_weight),
    .io_out_psum(PE_Array_6_20_io_out_psum)
  );
  basic_PE PE_Array_6_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_21_clock),
    .reset(PE_Array_6_21_reset),
    .io_in_activate(PE_Array_6_21_io_in_activate),
    .io_in_weight(PE_Array_6_21_io_in_weight),
    .io_in_psum(PE_Array_6_21_io_in_psum),
    .io_in_flow(PE_Array_6_21_io_in_flow),
    .io_in_shift(PE_Array_6_21_io_in_shift),
    .io_out_activate(PE_Array_6_21_io_out_activate),
    .io_out_weight(PE_Array_6_21_io_out_weight),
    .io_out_psum(PE_Array_6_21_io_out_psum)
  );
  basic_PE PE_Array_6_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_22_clock),
    .reset(PE_Array_6_22_reset),
    .io_in_activate(PE_Array_6_22_io_in_activate),
    .io_in_weight(PE_Array_6_22_io_in_weight),
    .io_in_psum(PE_Array_6_22_io_in_psum),
    .io_in_flow(PE_Array_6_22_io_in_flow),
    .io_in_shift(PE_Array_6_22_io_in_shift),
    .io_out_activate(PE_Array_6_22_io_out_activate),
    .io_out_weight(PE_Array_6_22_io_out_weight),
    .io_out_psum(PE_Array_6_22_io_out_psum)
  );
  basic_PE PE_Array_6_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_23_clock),
    .reset(PE_Array_6_23_reset),
    .io_in_activate(PE_Array_6_23_io_in_activate),
    .io_in_weight(PE_Array_6_23_io_in_weight),
    .io_in_psum(PE_Array_6_23_io_in_psum),
    .io_in_flow(PE_Array_6_23_io_in_flow),
    .io_in_shift(PE_Array_6_23_io_in_shift),
    .io_out_activate(PE_Array_6_23_io_out_activate),
    .io_out_weight(PE_Array_6_23_io_out_weight),
    .io_out_psum(PE_Array_6_23_io_out_psum)
  );
  basic_PE PE_Array_6_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_24_clock),
    .reset(PE_Array_6_24_reset),
    .io_in_activate(PE_Array_6_24_io_in_activate),
    .io_in_weight(PE_Array_6_24_io_in_weight),
    .io_in_psum(PE_Array_6_24_io_in_psum),
    .io_in_flow(PE_Array_6_24_io_in_flow),
    .io_in_shift(PE_Array_6_24_io_in_shift),
    .io_out_activate(PE_Array_6_24_io_out_activate),
    .io_out_weight(PE_Array_6_24_io_out_weight),
    .io_out_psum(PE_Array_6_24_io_out_psum)
  );
  basic_PE PE_Array_6_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_25_clock),
    .reset(PE_Array_6_25_reset),
    .io_in_activate(PE_Array_6_25_io_in_activate),
    .io_in_weight(PE_Array_6_25_io_in_weight),
    .io_in_psum(PE_Array_6_25_io_in_psum),
    .io_in_flow(PE_Array_6_25_io_in_flow),
    .io_in_shift(PE_Array_6_25_io_in_shift),
    .io_out_activate(PE_Array_6_25_io_out_activate),
    .io_out_weight(PE_Array_6_25_io_out_weight),
    .io_out_psum(PE_Array_6_25_io_out_psum)
  );
  basic_PE PE_Array_6_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_26_clock),
    .reset(PE_Array_6_26_reset),
    .io_in_activate(PE_Array_6_26_io_in_activate),
    .io_in_weight(PE_Array_6_26_io_in_weight),
    .io_in_psum(PE_Array_6_26_io_in_psum),
    .io_in_flow(PE_Array_6_26_io_in_flow),
    .io_in_shift(PE_Array_6_26_io_in_shift),
    .io_out_activate(PE_Array_6_26_io_out_activate),
    .io_out_weight(PE_Array_6_26_io_out_weight),
    .io_out_psum(PE_Array_6_26_io_out_psum)
  );
  basic_PE PE_Array_6_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_27_clock),
    .reset(PE_Array_6_27_reset),
    .io_in_activate(PE_Array_6_27_io_in_activate),
    .io_in_weight(PE_Array_6_27_io_in_weight),
    .io_in_psum(PE_Array_6_27_io_in_psum),
    .io_in_flow(PE_Array_6_27_io_in_flow),
    .io_in_shift(PE_Array_6_27_io_in_shift),
    .io_out_activate(PE_Array_6_27_io_out_activate),
    .io_out_weight(PE_Array_6_27_io_out_weight),
    .io_out_psum(PE_Array_6_27_io_out_psum)
  );
  basic_PE PE_Array_6_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_28_clock),
    .reset(PE_Array_6_28_reset),
    .io_in_activate(PE_Array_6_28_io_in_activate),
    .io_in_weight(PE_Array_6_28_io_in_weight),
    .io_in_psum(PE_Array_6_28_io_in_psum),
    .io_in_flow(PE_Array_6_28_io_in_flow),
    .io_in_shift(PE_Array_6_28_io_in_shift),
    .io_out_activate(PE_Array_6_28_io_out_activate),
    .io_out_weight(PE_Array_6_28_io_out_weight),
    .io_out_psum(PE_Array_6_28_io_out_psum)
  );
  basic_PE PE_Array_6_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_29_clock),
    .reset(PE_Array_6_29_reset),
    .io_in_activate(PE_Array_6_29_io_in_activate),
    .io_in_weight(PE_Array_6_29_io_in_weight),
    .io_in_psum(PE_Array_6_29_io_in_psum),
    .io_in_flow(PE_Array_6_29_io_in_flow),
    .io_in_shift(PE_Array_6_29_io_in_shift),
    .io_out_activate(PE_Array_6_29_io_out_activate),
    .io_out_weight(PE_Array_6_29_io_out_weight),
    .io_out_psum(PE_Array_6_29_io_out_psum)
  );
  basic_PE PE_Array_6_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_30_clock),
    .reset(PE_Array_6_30_reset),
    .io_in_activate(PE_Array_6_30_io_in_activate),
    .io_in_weight(PE_Array_6_30_io_in_weight),
    .io_in_psum(PE_Array_6_30_io_in_psum),
    .io_in_flow(PE_Array_6_30_io_in_flow),
    .io_in_shift(PE_Array_6_30_io_in_shift),
    .io_out_activate(PE_Array_6_30_io_out_activate),
    .io_out_weight(PE_Array_6_30_io_out_weight),
    .io_out_psum(PE_Array_6_30_io_out_psum)
  );
  basic_PE PE_Array_6_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_31_clock),
    .reset(PE_Array_6_31_reset),
    .io_in_activate(PE_Array_6_31_io_in_activate),
    .io_in_weight(PE_Array_6_31_io_in_weight),
    .io_in_psum(PE_Array_6_31_io_in_psum),
    .io_in_flow(PE_Array_6_31_io_in_flow),
    .io_in_shift(PE_Array_6_31_io_in_shift),
    .io_out_activate(PE_Array_6_31_io_out_activate),
    .io_out_weight(PE_Array_6_31_io_out_weight),
    .io_out_psum(PE_Array_6_31_io_out_psum)
  );
  basic_PE PE_Array_7_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_0_clock),
    .reset(PE_Array_7_0_reset),
    .io_in_activate(PE_Array_7_0_io_in_activate),
    .io_in_weight(PE_Array_7_0_io_in_weight),
    .io_in_psum(PE_Array_7_0_io_in_psum),
    .io_in_flow(PE_Array_7_0_io_in_flow),
    .io_in_shift(PE_Array_7_0_io_in_shift),
    .io_out_activate(PE_Array_7_0_io_out_activate),
    .io_out_weight(PE_Array_7_0_io_out_weight),
    .io_out_psum(PE_Array_7_0_io_out_psum)
  );
  basic_PE PE_Array_7_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_1_clock),
    .reset(PE_Array_7_1_reset),
    .io_in_activate(PE_Array_7_1_io_in_activate),
    .io_in_weight(PE_Array_7_1_io_in_weight),
    .io_in_psum(PE_Array_7_1_io_in_psum),
    .io_in_flow(PE_Array_7_1_io_in_flow),
    .io_in_shift(PE_Array_7_1_io_in_shift),
    .io_out_activate(PE_Array_7_1_io_out_activate),
    .io_out_weight(PE_Array_7_1_io_out_weight),
    .io_out_psum(PE_Array_7_1_io_out_psum)
  );
  basic_PE PE_Array_7_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_2_clock),
    .reset(PE_Array_7_2_reset),
    .io_in_activate(PE_Array_7_2_io_in_activate),
    .io_in_weight(PE_Array_7_2_io_in_weight),
    .io_in_psum(PE_Array_7_2_io_in_psum),
    .io_in_flow(PE_Array_7_2_io_in_flow),
    .io_in_shift(PE_Array_7_2_io_in_shift),
    .io_out_activate(PE_Array_7_2_io_out_activate),
    .io_out_weight(PE_Array_7_2_io_out_weight),
    .io_out_psum(PE_Array_7_2_io_out_psum)
  );
  basic_PE PE_Array_7_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_3_clock),
    .reset(PE_Array_7_3_reset),
    .io_in_activate(PE_Array_7_3_io_in_activate),
    .io_in_weight(PE_Array_7_3_io_in_weight),
    .io_in_psum(PE_Array_7_3_io_in_psum),
    .io_in_flow(PE_Array_7_3_io_in_flow),
    .io_in_shift(PE_Array_7_3_io_in_shift),
    .io_out_activate(PE_Array_7_3_io_out_activate),
    .io_out_weight(PE_Array_7_3_io_out_weight),
    .io_out_psum(PE_Array_7_3_io_out_psum)
  );
  basic_PE PE_Array_7_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_4_clock),
    .reset(PE_Array_7_4_reset),
    .io_in_activate(PE_Array_7_4_io_in_activate),
    .io_in_weight(PE_Array_7_4_io_in_weight),
    .io_in_psum(PE_Array_7_4_io_in_psum),
    .io_in_flow(PE_Array_7_4_io_in_flow),
    .io_in_shift(PE_Array_7_4_io_in_shift),
    .io_out_activate(PE_Array_7_4_io_out_activate),
    .io_out_weight(PE_Array_7_4_io_out_weight),
    .io_out_psum(PE_Array_7_4_io_out_psum)
  );
  basic_PE PE_Array_7_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_5_clock),
    .reset(PE_Array_7_5_reset),
    .io_in_activate(PE_Array_7_5_io_in_activate),
    .io_in_weight(PE_Array_7_5_io_in_weight),
    .io_in_psum(PE_Array_7_5_io_in_psum),
    .io_in_flow(PE_Array_7_5_io_in_flow),
    .io_in_shift(PE_Array_7_5_io_in_shift),
    .io_out_activate(PE_Array_7_5_io_out_activate),
    .io_out_weight(PE_Array_7_5_io_out_weight),
    .io_out_psum(PE_Array_7_5_io_out_psum)
  );
  basic_PE PE_Array_7_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_6_clock),
    .reset(PE_Array_7_6_reset),
    .io_in_activate(PE_Array_7_6_io_in_activate),
    .io_in_weight(PE_Array_7_6_io_in_weight),
    .io_in_psum(PE_Array_7_6_io_in_psum),
    .io_in_flow(PE_Array_7_6_io_in_flow),
    .io_in_shift(PE_Array_7_6_io_in_shift),
    .io_out_activate(PE_Array_7_6_io_out_activate),
    .io_out_weight(PE_Array_7_6_io_out_weight),
    .io_out_psum(PE_Array_7_6_io_out_psum)
  );
  basic_PE PE_Array_7_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_7_clock),
    .reset(PE_Array_7_7_reset),
    .io_in_activate(PE_Array_7_7_io_in_activate),
    .io_in_weight(PE_Array_7_7_io_in_weight),
    .io_in_psum(PE_Array_7_7_io_in_psum),
    .io_in_flow(PE_Array_7_7_io_in_flow),
    .io_in_shift(PE_Array_7_7_io_in_shift),
    .io_out_activate(PE_Array_7_7_io_out_activate),
    .io_out_weight(PE_Array_7_7_io_out_weight),
    .io_out_psum(PE_Array_7_7_io_out_psum)
  );
  basic_PE PE_Array_7_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_8_clock),
    .reset(PE_Array_7_8_reset),
    .io_in_activate(PE_Array_7_8_io_in_activate),
    .io_in_weight(PE_Array_7_8_io_in_weight),
    .io_in_psum(PE_Array_7_8_io_in_psum),
    .io_in_flow(PE_Array_7_8_io_in_flow),
    .io_in_shift(PE_Array_7_8_io_in_shift),
    .io_out_activate(PE_Array_7_8_io_out_activate),
    .io_out_weight(PE_Array_7_8_io_out_weight),
    .io_out_psum(PE_Array_7_8_io_out_psum)
  );
  basic_PE PE_Array_7_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_9_clock),
    .reset(PE_Array_7_9_reset),
    .io_in_activate(PE_Array_7_9_io_in_activate),
    .io_in_weight(PE_Array_7_9_io_in_weight),
    .io_in_psum(PE_Array_7_9_io_in_psum),
    .io_in_flow(PE_Array_7_9_io_in_flow),
    .io_in_shift(PE_Array_7_9_io_in_shift),
    .io_out_activate(PE_Array_7_9_io_out_activate),
    .io_out_weight(PE_Array_7_9_io_out_weight),
    .io_out_psum(PE_Array_7_9_io_out_psum)
  );
  basic_PE PE_Array_7_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_10_clock),
    .reset(PE_Array_7_10_reset),
    .io_in_activate(PE_Array_7_10_io_in_activate),
    .io_in_weight(PE_Array_7_10_io_in_weight),
    .io_in_psum(PE_Array_7_10_io_in_psum),
    .io_in_flow(PE_Array_7_10_io_in_flow),
    .io_in_shift(PE_Array_7_10_io_in_shift),
    .io_out_activate(PE_Array_7_10_io_out_activate),
    .io_out_weight(PE_Array_7_10_io_out_weight),
    .io_out_psum(PE_Array_7_10_io_out_psum)
  );
  basic_PE PE_Array_7_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_11_clock),
    .reset(PE_Array_7_11_reset),
    .io_in_activate(PE_Array_7_11_io_in_activate),
    .io_in_weight(PE_Array_7_11_io_in_weight),
    .io_in_psum(PE_Array_7_11_io_in_psum),
    .io_in_flow(PE_Array_7_11_io_in_flow),
    .io_in_shift(PE_Array_7_11_io_in_shift),
    .io_out_activate(PE_Array_7_11_io_out_activate),
    .io_out_weight(PE_Array_7_11_io_out_weight),
    .io_out_psum(PE_Array_7_11_io_out_psum)
  );
  basic_PE PE_Array_7_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_12_clock),
    .reset(PE_Array_7_12_reset),
    .io_in_activate(PE_Array_7_12_io_in_activate),
    .io_in_weight(PE_Array_7_12_io_in_weight),
    .io_in_psum(PE_Array_7_12_io_in_psum),
    .io_in_flow(PE_Array_7_12_io_in_flow),
    .io_in_shift(PE_Array_7_12_io_in_shift),
    .io_out_activate(PE_Array_7_12_io_out_activate),
    .io_out_weight(PE_Array_7_12_io_out_weight),
    .io_out_psum(PE_Array_7_12_io_out_psum)
  );
  basic_PE PE_Array_7_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_13_clock),
    .reset(PE_Array_7_13_reset),
    .io_in_activate(PE_Array_7_13_io_in_activate),
    .io_in_weight(PE_Array_7_13_io_in_weight),
    .io_in_psum(PE_Array_7_13_io_in_psum),
    .io_in_flow(PE_Array_7_13_io_in_flow),
    .io_in_shift(PE_Array_7_13_io_in_shift),
    .io_out_activate(PE_Array_7_13_io_out_activate),
    .io_out_weight(PE_Array_7_13_io_out_weight),
    .io_out_psum(PE_Array_7_13_io_out_psum)
  );
  basic_PE PE_Array_7_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_14_clock),
    .reset(PE_Array_7_14_reset),
    .io_in_activate(PE_Array_7_14_io_in_activate),
    .io_in_weight(PE_Array_7_14_io_in_weight),
    .io_in_psum(PE_Array_7_14_io_in_psum),
    .io_in_flow(PE_Array_7_14_io_in_flow),
    .io_in_shift(PE_Array_7_14_io_in_shift),
    .io_out_activate(PE_Array_7_14_io_out_activate),
    .io_out_weight(PE_Array_7_14_io_out_weight),
    .io_out_psum(PE_Array_7_14_io_out_psum)
  );
  basic_PE PE_Array_7_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_15_clock),
    .reset(PE_Array_7_15_reset),
    .io_in_activate(PE_Array_7_15_io_in_activate),
    .io_in_weight(PE_Array_7_15_io_in_weight),
    .io_in_psum(PE_Array_7_15_io_in_psum),
    .io_in_flow(PE_Array_7_15_io_in_flow),
    .io_in_shift(PE_Array_7_15_io_in_shift),
    .io_out_activate(PE_Array_7_15_io_out_activate),
    .io_out_weight(PE_Array_7_15_io_out_weight),
    .io_out_psum(PE_Array_7_15_io_out_psum)
  );
  basic_PE PE_Array_7_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_16_clock),
    .reset(PE_Array_7_16_reset),
    .io_in_activate(PE_Array_7_16_io_in_activate),
    .io_in_weight(PE_Array_7_16_io_in_weight),
    .io_in_psum(PE_Array_7_16_io_in_psum),
    .io_in_flow(PE_Array_7_16_io_in_flow),
    .io_in_shift(PE_Array_7_16_io_in_shift),
    .io_out_activate(PE_Array_7_16_io_out_activate),
    .io_out_weight(PE_Array_7_16_io_out_weight),
    .io_out_psum(PE_Array_7_16_io_out_psum)
  );
  basic_PE PE_Array_7_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_17_clock),
    .reset(PE_Array_7_17_reset),
    .io_in_activate(PE_Array_7_17_io_in_activate),
    .io_in_weight(PE_Array_7_17_io_in_weight),
    .io_in_psum(PE_Array_7_17_io_in_psum),
    .io_in_flow(PE_Array_7_17_io_in_flow),
    .io_in_shift(PE_Array_7_17_io_in_shift),
    .io_out_activate(PE_Array_7_17_io_out_activate),
    .io_out_weight(PE_Array_7_17_io_out_weight),
    .io_out_psum(PE_Array_7_17_io_out_psum)
  );
  basic_PE PE_Array_7_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_18_clock),
    .reset(PE_Array_7_18_reset),
    .io_in_activate(PE_Array_7_18_io_in_activate),
    .io_in_weight(PE_Array_7_18_io_in_weight),
    .io_in_psum(PE_Array_7_18_io_in_psum),
    .io_in_flow(PE_Array_7_18_io_in_flow),
    .io_in_shift(PE_Array_7_18_io_in_shift),
    .io_out_activate(PE_Array_7_18_io_out_activate),
    .io_out_weight(PE_Array_7_18_io_out_weight),
    .io_out_psum(PE_Array_7_18_io_out_psum)
  );
  basic_PE PE_Array_7_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_19_clock),
    .reset(PE_Array_7_19_reset),
    .io_in_activate(PE_Array_7_19_io_in_activate),
    .io_in_weight(PE_Array_7_19_io_in_weight),
    .io_in_psum(PE_Array_7_19_io_in_psum),
    .io_in_flow(PE_Array_7_19_io_in_flow),
    .io_in_shift(PE_Array_7_19_io_in_shift),
    .io_out_activate(PE_Array_7_19_io_out_activate),
    .io_out_weight(PE_Array_7_19_io_out_weight),
    .io_out_psum(PE_Array_7_19_io_out_psum)
  );
  basic_PE PE_Array_7_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_20_clock),
    .reset(PE_Array_7_20_reset),
    .io_in_activate(PE_Array_7_20_io_in_activate),
    .io_in_weight(PE_Array_7_20_io_in_weight),
    .io_in_psum(PE_Array_7_20_io_in_psum),
    .io_in_flow(PE_Array_7_20_io_in_flow),
    .io_in_shift(PE_Array_7_20_io_in_shift),
    .io_out_activate(PE_Array_7_20_io_out_activate),
    .io_out_weight(PE_Array_7_20_io_out_weight),
    .io_out_psum(PE_Array_7_20_io_out_psum)
  );
  basic_PE PE_Array_7_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_21_clock),
    .reset(PE_Array_7_21_reset),
    .io_in_activate(PE_Array_7_21_io_in_activate),
    .io_in_weight(PE_Array_7_21_io_in_weight),
    .io_in_psum(PE_Array_7_21_io_in_psum),
    .io_in_flow(PE_Array_7_21_io_in_flow),
    .io_in_shift(PE_Array_7_21_io_in_shift),
    .io_out_activate(PE_Array_7_21_io_out_activate),
    .io_out_weight(PE_Array_7_21_io_out_weight),
    .io_out_psum(PE_Array_7_21_io_out_psum)
  );
  basic_PE PE_Array_7_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_22_clock),
    .reset(PE_Array_7_22_reset),
    .io_in_activate(PE_Array_7_22_io_in_activate),
    .io_in_weight(PE_Array_7_22_io_in_weight),
    .io_in_psum(PE_Array_7_22_io_in_psum),
    .io_in_flow(PE_Array_7_22_io_in_flow),
    .io_in_shift(PE_Array_7_22_io_in_shift),
    .io_out_activate(PE_Array_7_22_io_out_activate),
    .io_out_weight(PE_Array_7_22_io_out_weight),
    .io_out_psum(PE_Array_7_22_io_out_psum)
  );
  basic_PE PE_Array_7_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_23_clock),
    .reset(PE_Array_7_23_reset),
    .io_in_activate(PE_Array_7_23_io_in_activate),
    .io_in_weight(PE_Array_7_23_io_in_weight),
    .io_in_psum(PE_Array_7_23_io_in_psum),
    .io_in_flow(PE_Array_7_23_io_in_flow),
    .io_in_shift(PE_Array_7_23_io_in_shift),
    .io_out_activate(PE_Array_7_23_io_out_activate),
    .io_out_weight(PE_Array_7_23_io_out_weight),
    .io_out_psum(PE_Array_7_23_io_out_psum)
  );
  basic_PE PE_Array_7_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_24_clock),
    .reset(PE_Array_7_24_reset),
    .io_in_activate(PE_Array_7_24_io_in_activate),
    .io_in_weight(PE_Array_7_24_io_in_weight),
    .io_in_psum(PE_Array_7_24_io_in_psum),
    .io_in_flow(PE_Array_7_24_io_in_flow),
    .io_in_shift(PE_Array_7_24_io_in_shift),
    .io_out_activate(PE_Array_7_24_io_out_activate),
    .io_out_weight(PE_Array_7_24_io_out_weight),
    .io_out_psum(PE_Array_7_24_io_out_psum)
  );
  basic_PE PE_Array_7_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_25_clock),
    .reset(PE_Array_7_25_reset),
    .io_in_activate(PE_Array_7_25_io_in_activate),
    .io_in_weight(PE_Array_7_25_io_in_weight),
    .io_in_psum(PE_Array_7_25_io_in_psum),
    .io_in_flow(PE_Array_7_25_io_in_flow),
    .io_in_shift(PE_Array_7_25_io_in_shift),
    .io_out_activate(PE_Array_7_25_io_out_activate),
    .io_out_weight(PE_Array_7_25_io_out_weight),
    .io_out_psum(PE_Array_7_25_io_out_psum)
  );
  basic_PE PE_Array_7_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_26_clock),
    .reset(PE_Array_7_26_reset),
    .io_in_activate(PE_Array_7_26_io_in_activate),
    .io_in_weight(PE_Array_7_26_io_in_weight),
    .io_in_psum(PE_Array_7_26_io_in_psum),
    .io_in_flow(PE_Array_7_26_io_in_flow),
    .io_in_shift(PE_Array_7_26_io_in_shift),
    .io_out_activate(PE_Array_7_26_io_out_activate),
    .io_out_weight(PE_Array_7_26_io_out_weight),
    .io_out_psum(PE_Array_7_26_io_out_psum)
  );
  basic_PE PE_Array_7_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_27_clock),
    .reset(PE_Array_7_27_reset),
    .io_in_activate(PE_Array_7_27_io_in_activate),
    .io_in_weight(PE_Array_7_27_io_in_weight),
    .io_in_psum(PE_Array_7_27_io_in_psum),
    .io_in_flow(PE_Array_7_27_io_in_flow),
    .io_in_shift(PE_Array_7_27_io_in_shift),
    .io_out_activate(PE_Array_7_27_io_out_activate),
    .io_out_weight(PE_Array_7_27_io_out_weight),
    .io_out_psum(PE_Array_7_27_io_out_psum)
  );
  basic_PE PE_Array_7_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_28_clock),
    .reset(PE_Array_7_28_reset),
    .io_in_activate(PE_Array_7_28_io_in_activate),
    .io_in_weight(PE_Array_7_28_io_in_weight),
    .io_in_psum(PE_Array_7_28_io_in_psum),
    .io_in_flow(PE_Array_7_28_io_in_flow),
    .io_in_shift(PE_Array_7_28_io_in_shift),
    .io_out_activate(PE_Array_7_28_io_out_activate),
    .io_out_weight(PE_Array_7_28_io_out_weight),
    .io_out_psum(PE_Array_7_28_io_out_psum)
  );
  basic_PE PE_Array_7_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_29_clock),
    .reset(PE_Array_7_29_reset),
    .io_in_activate(PE_Array_7_29_io_in_activate),
    .io_in_weight(PE_Array_7_29_io_in_weight),
    .io_in_psum(PE_Array_7_29_io_in_psum),
    .io_in_flow(PE_Array_7_29_io_in_flow),
    .io_in_shift(PE_Array_7_29_io_in_shift),
    .io_out_activate(PE_Array_7_29_io_out_activate),
    .io_out_weight(PE_Array_7_29_io_out_weight),
    .io_out_psum(PE_Array_7_29_io_out_psum)
  );
  basic_PE PE_Array_7_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_30_clock),
    .reset(PE_Array_7_30_reset),
    .io_in_activate(PE_Array_7_30_io_in_activate),
    .io_in_weight(PE_Array_7_30_io_in_weight),
    .io_in_psum(PE_Array_7_30_io_in_psum),
    .io_in_flow(PE_Array_7_30_io_in_flow),
    .io_in_shift(PE_Array_7_30_io_in_shift),
    .io_out_activate(PE_Array_7_30_io_out_activate),
    .io_out_weight(PE_Array_7_30_io_out_weight),
    .io_out_psum(PE_Array_7_30_io_out_psum)
  );
  basic_PE PE_Array_7_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_31_clock),
    .reset(PE_Array_7_31_reset),
    .io_in_activate(PE_Array_7_31_io_in_activate),
    .io_in_weight(PE_Array_7_31_io_in_weight),
    .io_in_psum(PE_Array_7_31_io_in_psum),
    .io_in_flow(PE_Array_7_31_io_in_flow),
    .io_in_shift(PE_Array_7_31_io_in_shift),
    .io_out_activate(PE_Array_7_31_io_out_activate),
    .io_out_weight(PE_Array_7_31_io_out_weight),
    .io_out_psum(PE_Array_7_31_io_out_psum)
  );
  basic_PE PE_Array_8_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_0_clock),
    .reset(PE_Array_8_0_reset),
    .io_in_activate(PE_Array_8_0_io_in_activate),
    .io_in_weight(PE_Array_8_0_io_in_weight),
    .io_in_psum(PE_Array_8_0_io_in_psum),
    .io_in_flow(PE_Array_8_0_io_in_flow),
    .io_in_shift(PE_Array_8_0_io_in_shift),
    .io_out_activate(PE_Array_8_0_io_out_activate),
    .io_out_weight(PE_Array_8_0_io_out_weight),
    .io_out_psum(PE_Array_8_0_io_out_psum)
  );
  basic_PE PE_Array_8_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_1_clock),
    .reset(PE_Array_8_1_reset),
    .io_in_activate(PE_Array_8_1_io_in_activate),
    .io_in_weight(PE_Array_8_1_io_in_weight),
    .io_in_psum(PE_Array_8_1_io_in_psum),
    .io_in_flow(PE_Array_8_1_io_in_flow),
    .io_in_shift(PE_Array_8_1_io_in_shift),
    .io_out_activate(PE_Array_8_1_io_out_activate),
    .io_out_weight(PE_Array_8_1_io_out_weight),
    .io_out_psum(PE_Array_8_1_io_out_psum)
  );
  basic_PE PE_Array_8_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_2_clock),
    .reset(PE_Array_8_2_reset),
    .io_in_activate(PE_Array_8_2_io_in_activate),
    .io_in_weight(PE_Array_8_2_io_in_weight),
    .io_in_psum(PE_Array_8_2_io_in_psum),
    .io_in_flow(PE_Array_8_2_io_in_flow),
    .io_in_shift(PE_Array_8_2_io_in_shift),
    .io_out_activate(PE_Array_8_2_io_out_activate),
    .io_out_weight(PE_Array_8_2_io_out_weight),
    .io_out_psum(PE_Array_8_2_io_out_psum)
  );
  basic_PE PE_Array_8_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_3_clock),
    .reset(PE_Array_8_3_reset),
    .io_in_activate(PE_Array_8_3_io_in_activate),
    .io_in_weight(PE_Array_8_3_io_in_weight),
    .io_in_psum(PE_Array_8_3_io_in_psum),
    .io_in_flow(PE_Array_8_3_io_in_flow),
    .io_in_shift(PE_Array_8_3_io_in_shift),
    .io_out_activate(PE_Array_8_3_io_out_activate),
    .io_out_weight(PE_Array_8_3_io_out_weight),
    .io_out_psum(PE_Array_8_3_io_out_psum)
  );
  basic_PE PE_Array_8_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_4_clock),
    .reset(PE_Array_8_4_reset),
    .io_in_activate(PE_Array_8_4_io_in_activate),
    .io_in_weight(PE_Array_8_4_io_in_weight),
    .io_in_psum(PE_Array_8_4_io_in_psum),
    .io_in_flow(PE_Array_8_4_io_in_flow),
    .io_in_shift(PE_Array_8_4_io_in_shift),
    .io_out_activate(PE_Array_8_4_io_out_activate),
    .io_out_weight(PE_Array_8_4_io_out_weight),
    .io_out_psum(PE_Array_8_4_io_out_psum)
  );
  basic_PE PE_Array_8_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_5_clock),
    .reset(PE_Array_8_5_reset),
    .io_in_activate(PE_Array_8_5_io_in_activate),
    .io_in_weight(PE_Array_8_5_io_in_weight),
    .io_in_psum(PE_Array_8_5_io_in_psum),
    .io_in_flow(PE_Array_8_5_io_in_flow),
    .io_in_shift(PE_Array_8_5_io_in_shift),
    .io_out_activate(PE_Array_8_5_io_out_activate),
    .io_out_weight(PE_Array_8_5_io_out_weight),
    .io_out_psum(PE_Array_8_5_io_out_psum)
  );
  basic_PE PE_Array_8_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_6_clock),
    .reset(PE_Array_8_6_reset),
    .io_in_activate(PE_Array_8_6_io_in_activate),
    .io_in_weight(PE_Array_8_6_io_in_weight),
    .io_in_psum(PE_Array_8_6_io_in_psum),
    .io_in_flow(PE_Array_8_6_io_in_flow),
    .io_in_shift(PE_Array_8_6_io_in_shift),
    .io_out_activate(PE_Array_8_6_io_out_activate),
    .io_out_weight(PE_Array_8_6_io_out_weight),
    .io_out_psum(PE_Array_8_6_io_out_psum)
  );
  basic_PE PE_Array_8_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_7_clock),
    .reset(PE_Array_8_7_reset),
    .io_in_activate(PE_Array_8_7_io_in_activate),
    .io_in_weight(PE_Array_8_7_io_in_weight),
    .io_in_psum(PE_Array_8_7_io_in_psum),
    .io_in_flow(PE_Array_8_7_io_in_flow),
    .io_in_shift(PE_Array_8_7_io_in_shift),
    .io_out_activate(PE_Array_8_7_io_out_activate),
    .io_out_weight(PE_Array_8_7_io_out_weight),
    .io_out_psum(PE_Array_8_7_io_out_psum)
  );
  basic_PE PE_Array_8_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_8_clock),
    .reset(PE_Array_8_8_reset),
    .io_in_activate(PE_Array_8_8_io_in_activate),
    .io_in_weight(PE_Array_8_8_io_in_weight),
    .io_in_psum(PE_Array_8_8_io_in_psum),
    .io_in_flow(PE_Array_8_8_io_in_flow),
    .io_in_shift(PE_Array_8_8_io_in_shift),
    .io_out_activate(PE_Array_8_8_io_out_activate),
    .io_out_weight(PE_Array_8_8_io_out_weight),
    .io_out_psum(PE_Array_8_8_io_out_psum)
  );
  basic_PE PE_Array_8_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_9_clock),
    .reset(PE_Array_8_9_reset),
    .io_in_activate(PE_Array_8_9_io_in_activate),
    .io_in_weight(PE_Array_8_9_io_in_weight),
    .io_in_psum(PE_Array_8_9_io_in_psum),
    .io_in_flow(PE_Array_8_9_io_in_flow),
    .io_in_shift(PE_Array_8_9_io_in_shift),
    .io_out_activate(PE_Array_8_9_io_out_activate),
    .io_out_weight(PE_Array_8_9_io_out_weight),
    .io_out_psum(PE_Array_8_9_io_out_psum)
  );
  basic_PE PE_Array_8_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_10_clock),
    .reset(PE_Array_8_10_reset),
    .io_in_activate(PE_Array_8_10_io_in_activate),
    .io_in_weight(PE_Array_8_10_io_in_weight),
    .io_in_psum(PE_Array_8_10_io_in_psum),
    .io_in_flow(PE_Array_8_10_io_in_flow),
    .io_in_shift(PE_Array_8_10_io_in_shift),
    .io_out_activate(PE_Array_8_10_io_out_activate),
    .io_out_weight(PE_Array_8_10_io_out_weight),
    .io_out_psum(PE_Array_8_10_io_out_psum)
  );
  basic_PE PE_Array_8_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_11_clock),
    .reset(PE_Array_8_11_reset),
    .io_in_activate(PE_Array_8_11_io_in_activate),
    .io_in_weight(PE_Array_8_11_io_in_weight),
    .io_in_psum(PE_Array_8_11_io_in_psum),
    .io_in_flow(PE_Array_8_11_io_in_flow),
    .io_in_shift(PE_Array_8_11_io_in_shift),
    .io_out_activate(PE_Array_8_11_io_out_activate),
    .io_out_weight(PE_Array_8_11_io_out_weight),
    .io_out_psum(PE_Array_8_11_io_out_psum)
  );
  basic_PE PE_Array_8_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_12_clock),
    .reset(PE_Array_8_12_reset),
    .io_in_activate(PE_Array_8_12_io_in_activate),
    .io_in_weight(PE_Array_8_12_io_in_weight),
    .io_in_psum(PE_Array_8_12_io_in_psum),
    .io_in_flow(PE_Array_8_12_io_in_flow),
    .io_in_shift(PE_Array_8_12_io_in_shift),
    .io_out_activate(PE_Array_8_12_io_out_activate),
    .io_out_weight(PE_Array_8_12_io_out_weight),
    .io_out_psum(PE_Array_8_12_io_out_psum)
  );
  basic_PE PE_Array_8_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_13_clock),
    .reset(PE_Array_8_13_reset),
    .io_in_activate(PE_Array_8_13_io_in_activate),
    .io_in_weight(PE_Array_8_13_io_in_weight),
    .io_in_psum(PE_Array_8_13_io_in_psum),
    .io_in_flow(PE_Array_8_13_io_in_flow),
    .io_in_shift(PE_Array_8_13_io_in_shift),
    .io_out_activate(PE_Array_8_13_io_out_activate),
    .io_out_weight(PE_Array_8_13_io_out_weight),
    .io_out_psum(PE_Array_8_13_io_out_psum)
  );
  basic_PE PE_Array_8_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_14_clock),
    .reset(PE_Array_8_14_reset),
    .io_in_activate(PE_Array_8_14_io_in_activate),
    .io_in_weight(PE_Array_8_14_io_in_weight),
    .io_in_psum(PE_Array_8_14_io_in_psum),
    .io_in_flow(PE_Array_8_14_io_in_flow),
    .io_in_shift(PE_Array_8_14_io_in_shift),
    .io_out_activate(PE_Array_8_14_io_out_activate),
    .io_out_weight(PE_Array_8_14_io_out_weight),
    .io_out_psum(PE_Array_8_14_io_out_psum)
  );
  basic_PE PE_Array_8_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_15_clock),
    .reset(PE_Array_8_15_reset),
    .io_in_activate(PE_Array_8_15_io_in_activate),
    .io_in_weight(PE_Array_8_15_io_in_weight),
    .io_in_psum(PE_Array_8_15_io_in_psum),
    .io_in_flow(PE_Array_8_15_io_in_flow),
    .io_in_shift(PE_Array_8_15_io_in_shift),
    .io_out_activate(PE_Array_8_15_io_out_activate),
    .io_out_weight(PE_Array_8_15_io_out_weight),
    .io_out_psum(PE_Array_8_15_io_out_psum)
  );
  basic_PE PE_Array_8_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_16_clock),
    .reset(PE_Array_8_16_reset),
    .io_in_activate(PE_Array_8_16_io_in_activate),
    .io_in_weight(PE_Array_8_16_io_in_weight),
    .io_in_psum(PE_Array_8_16_io_in_psum),
    .io_in_flow(PE_Array_8_16_io_in_flow),
    .io_in_shift(PE_Array_8_16_io_in_shift),
    .io_out_activate(PE_Array_8_16_io_out_activate),
    .io_out_weight(PE_Array_8_16_io_out_weight),
    .io_out_psum(PE_Array_8_16_io_out_psum)
  );
  basic_PE PE_Array_8_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_17_clock),
    .reset(PE_Array_8_17_reset),
    .io_in_activate(PE_Array_8_17_io_in_activate),
    .io_in_weight(PE_Array_8_17_io_in_weight),
    .io_in_psum(PE_Array_8_17_io_in_psum),
    .io_in_flow(PE_Array_8_17_io_in_flow),
    .io_in_shift(PE_Array_8_17_io_in_shift),
    .io_out_activate(PE_Array_8_17_io_out_activate),
    .io_out_weight(PE_Array_8_17_io_out_weight),
    .io_out_psum(PE_Array_8_17_io_out_psum)
  );
  basic_PE PE_Array_8_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_18_clock),
    .reset(PE_Array_8_18_reset),
    .io_in_activate(PE_Array_8_18_io_in_activate),
    .io_in_weight(PE_Array_8_18_io_in_weight),
    .io_in_psum(PE_Array_8_18_io_in_psum),
    .io_in_flow(PE_Array_8_18_io_in_flow),
    .io_in_shift(PE_Array_8_18_io_in_shift),
    .io_out_activate(PE_Array_8_18_io_out_activate),
    .io_out_weight(PE_Array_8_18_io_out_weight),
    .io_out_psum(PE_Array_8_18_io_out_psum)
  );
  basic_PE PE_Array_8_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_19_clock),
    .reset(PE_Array_8_19_reset),
    .io_in_activate(PE_Array_8_19_io_in_activate),
    .io_in_weight(PE_Array_8_19_io_in_weight),
    .io_in_psum(PE_Array_8_19_io_in_psum),
    .io_in_flow(PE_Array_8_19_io_in_flow),
    .io_in_shift(PE_Array_8_19_io_in_shift),
    .io_out_activate(PE_Array_8_19_io_out_activate),
    .io_out_weight(PE_Array_8_19_io_out_weight),
    .io_out_psum(PE_Array_8_19_io_out_psum)
  );
  basic_PE PE_Array_8_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_20_clock),
    .reset(PE_Array_8_20_reset),
    .io_in_activate(PE_Array_8_20_io_in_activate),
    .io_in_weight(PE_Array_8_20_io_in_weight),
    .io_in_psum(PE_Array_8_20_io_in_psum),
    .io_in_flow(PE_Array_8_20_io_in_flow),
    .io_in_shift(PE_Array_8_20_io_in_shift),
    .io_out_activate(PE_Array_8_20_io_out_activate),
    .io_out_weight(PE_Array_8_20_io_out_weight),
    .io_out_psum(PE_Array_8_20_io_out_psum)
  );
  basic_PE PE_Array_8_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_21_clock),
    .reset(PE_Array_8_21_reset),
    .io_in_activate(PE_Array_8_21_io_in_activate),
    .io_in_weight(PE_Array_8_21_io_in_weight),
    .io_in_psum(PE_Array_8_21_io_in_psum),
    .io_in_flow(PE_Array_8_21_io_in_flow),
    .io_in_shift(PE_Array_8_21_io_in_shift),
    .io_out_activate(PE_Array_8_21_io_out_activate),
    .io_out_weight(PE_Array_8_21_io_out_weight),
    .io_out_psum(PE_Array_8_21_io_out_psum)
  );
  basic_PE PE_Array_8_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_22_clock),
    .reset(PE_Array_8_22_reset),
    .io_in_activate(PE_Array_8_22_io_in_activate),
    .io_in_weight(PE_Array_8_22_io_in_weight),
    .io_in_psum(PE_Array_8_22_io_in_psum),
    .io_in_flow(PE_Array_8_22_io_in_flow),
    .io_in_shift(PE_Array_8_22_io_in_shift),
    .io_out_activate(PE_Array_8_22_io_out_activate),
    .io_out_weight(PE_Array_8_22_io_out_weight),
    .io_out_psum(PE_Array_8_22_io_out_psum)
  );
  basic_PE PE_Array_8_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_23_clock),
    .reset(PE_Array_8_23_reset),
    .io_in_activate(PE_Array_8_23_io_in_activate),
    .io_in_weight(PE_Array_8_23_io_in_weight),
    .io_in_psum(PE_Array_8_23_io_in_psum),
    .io_in_flow(PE_Array_8_23_io_in_flow),
    .io_in_shift(PE_Array_8_23_io_in_shift),
    .io_out_activate(PE_Array_8_23_io_out_activate),
    .io_out_weight(PE_Array_8_23_io_out_weight),
    .io_out_psum(PE_Array_8_23_io_out_psum)
  );
  basic_PE PE_Array_8_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_24_clock),
    .reset(PE_Array_8_24_reset),
    .io_in_activate(PE_Array_8_24_io_in_activate),
    .io_in_weight(PE_Array_8_24_io_in_weight),
    .io_in_psum(PE_Array_8_24_io_in_psum),
    .io_in_flow(PE_Array_8_24_io_in_flow),
    .io_in_shift(PE_Array_8_24_io_in_shift),
    .io_out_activate(PE_Array_8_24_io_out_activate),
    .io_out_weight(PE_Array_8_24_io_out_weight),
    .io_out_psum(PE_Array_8_24_io_out_psum)
  );
  basic_PE PE_Array_8_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_25_clock),
    .reset(PE_Array_8_25_reset),
    .io_in_activate(PE_Array_8_25_io_in_activate),
    .io_in_weight(PE_Array_8_25_io_in_weight),
    .io_in_psum(PE_Array_8_25_io_in_psum),
    .io_in_flow(PE_Array_8_25_io_in_flow),
    .io_in_shift(PE_Array_8_25_io_in_shift),
    .io_out_activate(PE_Array_8_25_io_out_activate),
    .io_out_weight(PE_Array_8_25_io_out_weight),
    .io_out_psum(PE_Array_8_25_io_out_psum)
  );
  basic_PE PE_Array_8_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_26_clock),
    .reset(PE_Array_8_26_reset),
    .io_in_activate(PE_Array_8_26_io_in_activate),
    .io_in_weight(PE_Array_8_26_io_in_weight),
    .io_in_psum(PE_Array_8_26_io_in_psum),
    .io_in_flow(PE_Array_8_26_io_in_flow),
    .io_in_shift(PE_Array_8_26_io_in_shift),
    .io_out_activate(PE_Array_8_26_io_out_activate),
    .io_out_weight(PE_Array_8_26_io_out_weight),
    .io_out_psum(PE_Array_8_26_io_out_psum)
  );
  basic_PE PE_Array_8_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_27_clock),
    .reset(PE_Array_8_27_reset),
    .io_in_activate(PE_Array_8_27_io_in_activate),
    .io_in_weight(PE_Array_8_27_io_in_weight),
    .io_in_psum(PE_Array_8_27_io_in_psum),
    .io_in_flow(PE_Array_8_27_io_in_flow),
    .io_in_shift(PE_Array_8_27_io_in_shift),
    .io_out_activate(PE_Array_8_27_io_out_activate),
    .io_out_weight(PE_Array_8_27_io_out_weight),
    .io_out_psum(PE_Array_8_27_io_out_psum)
  );
  basic_PE PE_Array_8_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_28_clock),
    .reset(PE_Array_8_28_reset),
    .io_in_activate(PE_Array_8_28_io_in_activate),
    .io_in_weight(PE_Array_8_28_io_in_weight),
    .io_in_psum(PE_Array_8_28_io_in_psum),
    .io_in_flow(PE_Array_8_28_io_in_flow),
    .io_in_shift(PE_Array_8_28_io_in_shift),
    .io_out_activate(PE_Array_8_28_io_out_activate),
    .io_out_weight(PE_Array_8_28_io_out_weight),
    .io_out_psum(PE_Array_8_28_io_out_psum)
  );
  basic_PE PE_Array_8_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_29_clock),
    .reset(PE_Array_8_29_reset),
    .io_in_activate(PE_Array_8_29_io_in_activate),
    .io_in_weight(PE_Array_8_29_io_in_weight),
    .io_in_psum(PE_Array_8_29_io_in_psum),
    .io_in_flow(PE_Array_8_29_io_in_flow),
    .io_in_shift(PE_Array_8_29_io_in_shift),
    .io_out_activate(PE_Array_8_29_io_out_activate),
    .io_out_weight(PE_Array_8_29_io_out_weight),
    .io_out_psum(PE_Array_8_29_io_out_psum)
  );
  basic_PE PE_Array_8_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_30_clock),
    .reset(PE_Array_8_30_reset),
    .io_in_activate(PE_Array_8_30_io_in_activate),
    .io_in_weight(PE_Array_8_30_io_in_weight),
    .io_in_psum(PE_Array_8_30_io_in_psum),
    .io_in_flow(PE_Array_8_30_io_in_flow),
    .io_in_shift(PE_Array_8_30_io_in_shift),
    .io_out_activate(PE_Array_8_30_io_out_activate),
    .io_out_weight(PE_Array_8_30_io_out_weight),
    .io_out_psum(PE_Array_8_30_io_out_psum)
  );
  basic_PE PE_Array_8_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_8_31_clock),
    .reset(PE_Array_8_31_reset),
    .io_in_activate(PE_Array_8_31_io_in_activate),
    .io_in_weight(PE_Array_8_31_io_in_weight),
    .io_in_psum(PE_Array_8_31_io_in_psum),
    .io_in_flow(PE_Array_8_31_io_in_flow),
    .io_in_shift(PE_Array_8_31_io_in_shift),
    .io_out_activate(PE_Array_8_31_io_out_activate),
    .io_out_weight(PE_Array_8_31_io_out_weight),
    .io_out_psum(PE_Array_8_31_io_out_psum)
  );
  basic_PE PE_Array_9_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_0_clock),
    .reset(PE_Array_9_0_reset),
    .io_in_activate(PE_Array_9_0_io_in_activate),
    .io_in_weight(PE_Array_9_0_io_in_weight),
    .io_in_psum(PE_Array_9_0_io_in_psum),
    .io_in_flow(PE_Array_9_0_io_in_flow),
    .io_in_shift(PE_Array_9_0_io_in_shift),
    .io_out_activate(PE_Array_9_0_io_out_activate),
    .io_out_weight(PE_Array_9_0_io_out_weight),
    .io_out_psum(PE_Array_9_0_io_out_psum)
  );
  basic_PE PE_Array_9_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_1_clock),
    .reset(PE_Array_9_1_reset),
    .io_in_activate(PE_Array_9_1_io_in_activate),
    .io_in_weight(PE_Array_9_1_io_in_weight),
    .io_in_psum(PE_Array_9_1_io_in_psum),
    .io_in_flow(PE_Array_9_1_io_in_flow),
    .io_in_shift(PE_Array_9_1_io_in_shift),
    .io_out_activate(PE_Array_9_1_io_out_activate),
    .io_out_weight(PE_Array_9_1_io_out_weight),
    .io_out_psum(PE_Array_9_1_io_out_psum)
  );
  basic_PE PE_Array_9_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_2_clock),
    .reset(PE_Array_9_2_reset),
    .io_in_activate(PE_Array_9_2_io_in_activate),
    .io_in_weight(PE_Array_9_2_io_in_weight),
    .io_in_psum(PE_Array_9_2_io_in_psum),
    .io_in_flow(PE_Array_9_2_io_in_flow),
    .io_in_shift(PE_Array_9_2_io_in_shift),
    .io_out_activate(PE_Array_9_2_io_out_activate),
    .io_out_weight(PE_Array_9_2_io_out_weight),
    .io_out_psum(PE_Array_9_2_io_out_psum)
  );
  basic_PE PE_Array_9_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_3_clock),
    .reset(PE_Array_9_3_reset),
    .io_in_activate(PE_Array_9_3_io_in_activate),
    .io_in_weight(PE_Array_9_3_io_in_weight),
    .io_in_psum(PE_Array_9_3_io_in_psum),
    .io_in_flow(PE_Array_9_3_io_in_flow),
    .io_in_shift(PE_Array_9_3_io_in_shift),
    .io_out_activate(PE_Array_9_3_io_out_activate),
    .io_out_weight(PE_Array_9_3_io_out_weight),
    .io_out_psum(PE_Array_9_3_io_out_psum)
  );
  basic_PE PE_Array_9_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_4_clock),
    .reset(PE_Array_9_4_reset),
    .io_in_activate(PE_Array_9_4_io_in_activate),
    .io_in_weight(PE_Array_9_4_io_in_weight),
    .io_in_psum(PE_Array_9_4_io_in_psum),
    .io_in_flow(PE_Array_9_4_io_in_flow),
    .io_in_shift(PE_Array_9_4_io_in_shift),
    .io_out_activate(PE_Array_9_4_io_out_activate),
    .io_out_weight(PE_Array_9_4_io_out_weight),
    .io_out_psum(PE_Array_9_4_io_out_psum)
  );
  basic_PE PE_Array_9_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_5_clock),
    .reset(PE_Array_9_5_reset),
    .io_in_activate(PE_Array_9_5_io_in_activate),
    .io_in_weight(PE_Array_9_5_io_in_weight),
    .io_in_psum(PE_Array_9_5_io_in_psum),
    .io_in_flow(PE_Array_9_5_io_in_flow),
    .io_in_shift(PE_Array_9_5_io_in_shift),
    .io_out_activate(PE_Array_9_5_io_out_activate),
    .io_out_weight(PE_Array_9_5_io_out_weight),
    .io_out_psum(PE_Array_9_5_io_out_psum)
  );
  basic_PE PE_Array_9_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_6_clock),
    .reset(PE_Array_9_6_reset),
    .io_in_activate(PE_Array_9_6_io_in_activate),
    .io_in_weight(PE_Array_9_6_io_in_weight),
    .io_in_psum(PE_Array_9_6_io_in_psum),
    .io_in_flow(PE_Array_9_6_io_in_flow),
    .io_in_shift(PE_Array_9_6_io_in_shift),
    .io_out_activate(PE_Array_9_6_io_out_activate),
    .io_out_weight(PE_Array_9_6_io_out_weight),
    .io_out_psum(PE_Array_9_6_io_out_psum)
  );
  basic_PE PE_Array_9_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_7_clock),
    .reset(PE_Array_9_7_reset),
    .io_in_activate(PE_Array_9_7_io_in_activate),
    .io_in_weight(PE_Array_9_7_io_in_weight),
    .io_in_psum(PE_Array_9_7_io_in_psum),
    .io_in_flow(PE_Array_9_7_io_in_flow),
    .io_in_shift(PE_Array_9_7_io_in_shift),
    .io_out_activate(PE_Array_9_7_io_out_activate),
    .io_out_weight(PE_Array_9_7_io_out_weight),
    .io_out_psum(PE_Array_9_7_io_out_psum)
  );
  basic_PE PE_Array_9_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_8_clock),
    .reset(PE_Array_9_8_reset),
    .io_in_activate(PE_Array_9_8_io_in_activate),
    .io_in_weight(PE_Array_9_8_io_in_weight),
    .io_in_psum(PE_Array_9_8_io_in_psum),
    .io_in_flow(PE_Array_9_8_io_in_flow),
    .io_in_shift(PE_Array_9_8_io_in_shift),
    .io_out_activate(PE_Array_9_8_io_out_activate),
    .io_out_weight(PE_Array_9_8_io_out_weight),
    .io_out_psum(PE_Array_9_8_io_out_psum)
  );
  basic_PE PE_Array_9_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_9_clock),
    .reset(PE_Array_9_9_reset),
    .io_in_activate(PE_Array_9_9_io_in_activate),
    .io_in_weight(PE_Array_9_9_io_in_weight),
    .io_in_psum(PE_Array_9_9_io_in_psum),
    .io_in_flow(PE_Array_9_9_io_in_flow),
    .io_in_shift(PE_Array_9_9_io_in_shift),
    .io_out_activate(PE_Array_9_9_io_out_activate),
    .io_out_weight(PE_Array_9_9_io_out_weight),
    .io_out_psum(PE_Array_9_9_io_out_psum)
  );
  basic_PE PE_Array_9_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_10_clock),
    .reset(PE_Array_9_10_reset),
    .io_in_activate(PE_Array_9_10_io_in_activate),
    .io_in_weight(PE_Array_9_10_io_in_weight),
    .io_in_psum(PE_Array_9_10_io_in_psum),
    .io_in_flow(PE_Array_9_10_io_in_flow),
    .io_in_shift(PE_Array_9_10_io_in_shift),
    .io_out_activate(PE_Array_9_10_io_out_activate),
    .io_out_weight(PE_Array_9_10_io_out_weight),
    .io_out_psum(PE_Array_9_10_io_out_psum)
  );
  basic_PE PE_Array_9_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_11_clock),
    .reset(PE_Array_9_11_reset),
    .io_in_activate(PE_Array_9_11_io_in_activate),
    .io_in_weight(PE_Array_9_11_io_in_weight),
    .io_in_psum(PE_Array_9_11_io_in_psum),
    .io_in_flow(PE_Array_9_11_io_in_flow),
    .io_in_shift(PE_Array_9_11_io_in_shift),
    .io_out_activate(PE_Array_9_11_io_out_activate),
    .io_out_weight(PE_Array_9_11_io_out_weight),
    .io_out_psum(PE_Array_9_11_io_out_psum)
  );
  basic_PE PE_Array_9_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_12_clock),
    .reset(PE_Array_9_12_reset),
    .io_in_activate(PE_Array_9_12_io_in_activate),
    .io_in_weight(PE_Array_9_12_io_in_weight),
    .io_in_psum(PE_Array_9_12_io_in_psum),
    .io_in_flow(PE_Array_9_12_io_in_flow),
    .io_in_shift(PE_Array_9_12_io_in_shift),
    .io_out_activate(PE_Array_9_12_io_out_activate),
    .io_out_weight(PE_Array_9_12_io_out_weight),
    .io_out_psum(PE_Array_9_12_io_out_psum)
  );
  basic_PE PE_Array_9_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_13_clock),
    .reset(PE_Array_9_13_reset),
    .io_in_activate(PE_Array_9_13_io_in_activate),
    .io_in_weight(PE_Array_9_13_io_in_weight),
    .io_in_psum(PE_Array_9_13_io_in_psum),
    .io_in_flow(PE_Array_9_13_io_in_flow),
    .io_in_shift(PE_Array_9_13_io_in_shift),
    .io_out_activate(PE_Array_9_13_io_out_activate),
    .io_out_weight(PE_Array_9_13_io_out_weight),
    .io_out_psum(PE_Array_9_13_io_out_psum)
  );
  basic_PE PE_Array_9_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_14_clock),
    .reset(PE_Array_9_14_reset),
    .io_in_activate(PE_Array_9_14_io_in_activate),
    .io_in_weight(PE_Array_9_14_io_in_weight),
    .io_in_psum(PE_Array_9_14_io_in_psum),
    .io_in_flow(PE_Array_9_14_io_in_flow),
    .io_in_shift(PE_Array_9_14_io_in_shift),
    .io_out_activate(PE_Array_9_14_io_out_activate),
    .io_out_weight(PE_Array_9_14_io_out_weight),
    .io_out_psum(PE_Array_9_14_io_out_psum)
  );
  basic_PE PE_Array_9_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_15_clock),
    .reset(PE_Array_9_15_reset),
    .io_in_activate(PE_Array_9_15_io_in_activate),
    .io_in_weight(PE_Array_9_15_io_in_weight),
    .io_in_psum(PE_Array_9_15_io_in_psum),
    .io_in_flow(PE_Array_9_15_io_in_flow),
    .io_in_shift(PE_Array_9_15_io_in_shift),
    .io_out_activate(PE_Array_9_15_io_out_activate),
    .io_out_weight(PE_Array_9_15_io_out_weight),
    .io_out_psum(PE_Array_9_15_io_out_psum)
  );
  basic_PE PE_Array_9_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_16_clock),
    .reset(PE_Array_9_16_reset),
    .io_in_activate(PE_Array_9_16_io_in_activate),
    .io_in_weight(PE_Array_9_16_io_in_weight),
    .io_in_psum(PE_Array_9_16_io_in_psum),
    .io_in_flow(PE_Array_9_16_io_in_flow),
    .io_in_shift(PE_Array_9_16_io_in_shift),
    .io_out_activate(PE_Array_9_16_io_out_activate),
    .io_out_weight(PE_Array_9_16_io_out_weight),
    .io_out_psum(PE_Array_9_16_io_out_psum)
  );
  basic_PE PE_Array_9_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_17_clock),
    .reset(PE_Array_9_17_reset),
    .io_in_activate(PE_Array_9_17_io_in_activate),
    .io_in_weight(PE_Array_9_17_io_in_weight),
    .io_in_psum(PE_Array_9_17_io_in_psum),
    .io_in_flow(PE_Array_9_17_io_in_flow),
    .io_in_shift(PE_Array_9_17_io_in_shift),
    .io_out_activate(PE_Array_9_17_io_out_activate),
    .io_out_weight(PE_Array_9_17_io_out_weight),
    .io_out_psum(PE_Array_9_17_io_out_psum)
  );
  basic_PE PE_Array_9_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_18_clock),
    .reset(PE_Array_9_18_reset),
    .io_in_activate(PE_Array_9_18_io_in_activate),
    .io_in_weight(PE_Array_9_18_io_in_weight),
    .io_in_psum(PE_Array_9_18_io_in_psum),
    .io_in_flow(PE_Array_9_18_io_in_flow),
    .io_in_shift(PE_Array_9_18_io_in_shift),
    .io_out_activate(PE_Array_9_18_io_out_activate),
    .io_out_weight(PE_Array_9_18_io_out_weight),
    .io_out_psum(PE_Array_9_18_io_out_psum)
  );
  basic_PE PE_Array_9_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_19_clock),
    .reset(PE_Array_9_19_reset),
    .io_in_activate(PE_Array_9_19_io_in_activate),
    .io_in_weight(PE_Array_9_19_io_in_weight),
    .io_in_psum(PE_Array_9_19_io_in_psum),
    .io_in_flow(PE_Array_9_19_io_in_flow),
    .io_in_shift(PE_Array_9_19_io_in_shift),
    .io_out_activate(PE_Array_9_19_io_out_activate),
    .io_out_weight(PE_Array_9_19_io_out_weight),
    .io_out_psum(PE_Array_9_19_io_out_psum)
  );
  basic_PE PE_Array_9_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_20_clock),
    .reset(PE_Array_9_20_reset),
    .io_in_activate(PE_Array_9_20_io_in_activate),
    .io_in_weight(PE_Array_9_20_io_in_weight),
    .io_in_psum(PE_Array_9_20_io_in_psum),
    .io_in_flow(PE_Array_9_20_io_in_flow),
    .io_in_shift(PE_Array_9_20_io_in_shift),
    .io_out_activate(PE_Array_9_20_io_out_activate),
    .io_out_weight(PE_Array_9_20_io_out_weight),
    .io_out_psum(PE_Array_9_20_io_out_psum)
  );
  basic_PE PE_Array_9_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_21_clock),
    .reset(PE_Array_9_21_reset),
    .io_in_activate(PE_Array_9_21_io_in_activate),
    .io_in_weight(PE_Array_9_21_io_in_weight),
    .io_in_psum(PE_Array_9_21_io_in_psum),
    .io_in_flow(PE_Array_9_21_io_in_flow),
    .io_in_shift(PE_Array_9_21_io_in_shift),
    .io_out_activate(PE_Array_9_21_io_out_activate),
    .io_out_weight(PE_Array_9_21_io_out_weight),
    .io_out_psum(PE_Array_9_21_io_out_psum)
  );
  basic_PE PE_Array_9_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_22_clock),
    .reset(PE_Array_9_22_reset),
    .io_in_activate(PE_Array_9_22_io_in_activate),
    .io_in_weight(PE_Array_9_22_io_in_weight),
    .io_in_psum(PE_Array_9_22_io_in_psum),
    .io_in_flow(PE_Array_9_22_io_in_flow),
    .io_in_shift(PE_Array_9_22_io_in_shift),
    .io_out_activate(PE_Array_9_22_io_out_activate),
    .io_out_weight(PE_Array_9_22_io_out_weight),
    .io_out_psum(PE_Array_9_22_io_out_psum)
  );
  basic_PE PE_Array_9_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_23_clock),
    .reset(PE_Array_9_23_reset),
    .io_in_activate(PE_Array_9_23_io_in_activate),
    .io_in_weight(PE_Array_9_23_io_in_weight),
    .io_in_psum(PE_Array_9_23_io_in_psum),
    .io_in_flow(PE_Array_9_23_io_in_flow),
    .io_in_shift(PE_Array_9_23_io_in_shift),
    .io_out_activate(PE_Array_9_23_io_out_activate),
    .io_out_weight(PE_Array_9_23_io_out_weight),
    .io_out_psum(PE_Array_9_23_io_out_psum)
  );
  basic_PE PE_Array_9_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_24_clock),
    .reset(PE_Array_9_24_reset),
    .io_in_activate(PE_Array_9_24_io_in_activate),
    .io_in_weight(PE_Array_9_24_io_in_weight),
    .io_in_psum(PE_Array_9_24_io_in_psum),
    .io_in_flow(PE_Array_9_24_io_in_flow),
    .io_in_shift(PE_Array_9_24_io_in_shift),
    .io_out_activate(PE_Array_9_24_io_out_activate),
    .io_out_weight(PE_Array_9_24_io_out_weight),
    .io_out_psum(PE_Array_9_24_io_out_psum)
  );
  basic_PE PE_Array_9_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_25_clock),
    .reset(PE_Array_9_25_reset),
    .io_in_activate(PE_Array_9_25_io_in_activate),
    .io_in_weight(PE_Array_9_25_io_in_weight),
    .io_in_psum(PE_Array_9_25_io_in_psum),
    .io_in_flow(PE_Array_9_25_io_in_flow),
    .io_in_shift(PE_Array_9_25_io_in_shift),
    .io_out_activate(PE_Array_9_25_io_out_activate),
    .io_out_weight(PE_Array_9_25_io_out_weight),
    .io_out_psum(PE_Array_9_25_io_out_psum)
  );
  basic_PE PE_Array_9_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_26_clock),
    .reset(PE_Array_9_26_reset),
    .io_in_activate(PE_Array_9_26_io_in_activate),
    .io_in_weight(PE_Array_9_26_io_in_weight),
    .io_in_psum(PE_Array_9_26_io_in_psum),
    .io_in_flow(PE_Array_9_26_io_in_flow),
    .io_in_shift(PE_Array_9_26_io_in_shift),
    .io_out_activate(PE_Array_9_26_io_out_activate),
    .io_out_weight(PE_Array_9_26_io_out_weight),
    .io_out_psum(PE_Array_9_26_io_out_psum)
  );
  basic_PE PE_Array_9_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_27_clock),
    .reset(PE_Array_9_27_reset),
    .io_in_activate(PE_Array_9_27_io_in_activate),
    .io_in_weight(PE_Array_9_27_io_in_weight),
    .io_in_psum(PE_Array_9_27_io_in_psum),
    .io_in_flow(PE_Array_9_27_io_in_flow),
    .io_in_shift(PE_Array_9_27_io_in_shift),
    .io_out_activate(PE_Array_9_27_io_out_activate),
    .io_out_weight(PE_Array_9_27_io_out_weight),
    .io_out_psum(PE_Array_9_27_io_out_psum)
  );
  basic_PE PE_Array_9_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_28_clock),
    .reset(PE_Array_9_28_reset),
    .io_in_activate(PE_Array_9_28_io_in_activate),
    .io_in_weight(PE_Array_9_28_io_in_weight),
    .io_in_psum(PE_Array_9_28_io_in_psum),
    .io_in_flow(PE_Array_9_28_io_in_flow),
    .io_in_shift(PE_Array_9_28_io_in_shift),
    .io_out_activate(PE_Array_9_28_io_out_activate),
    .io_out_weight(PE_Array_9_28_io_out_weight),
    .io_out_psum(PE_Array_9_28_io_out_psum)
  );
  basic_PE PE_Array_9_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_29_clock),
    .reset(PE_Array_9_29_reset),
    .io_in_activate(PE_Array_9_29_io_in_activate),
    .io_in_weight(PE_Array_9_29_io_in_weight),
    .io_in_psum(PE_Array_9_29_io_in_psum),
    .io_in_flow(PE_Array_9_29_io_in_flow),
    .io_in_shift(PE_Array_9_29_io_in_shift),
    .io_out_activate(PE_Array_9_29_io_out_activate),
    .io_out_weight(PE_Array_9_29_io_out_weight),
    .io_out_psum(PE_Array_9_29_io_out_psum)
  );
  basic_PE PE_Array_9_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_30_clock),
    .reset(PE_Array_9_30_reset),
    .io_in_activate(PE_Array_9_30_io_in_activate),
    .io_in_weight(PE_Array_9_30_io_in_weight),
    .io_in_psum(PE_Array_9_30_io_in_psum),
    .io_in_flow(PE_Array_9_30_io_in_flow),
    .io_in_shift(PE_Array_9_30_io_in_shift),
    .io_out_activate(PE_Array_9_30_io_out_activate),
    .io_out_weight(PE_Array_9_30_io_out_weight),
    .io_out_psum(PE_Array_9_30_io_out_psum)
  );
  basic_PE PE_Array_9_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_9_31_clock),
    .reset(PE_Array_9_31_reset),
    .io_in_activate(PE_Array_9_31_io_in_activate),
    .io_in_weight(PE_Array_9_31_io_in_weight),
    .io_in_psum(PE_Array_9_31_io_in_psum),
    .io_in_flow(PE_Array_9_31_io_in_flow),
    .io_in_shift(PE_Array_9_31_io_in_shift),
    .io_out_activate(PE_Array_9_31_io_out_activate),
    .io_out_weight(PE_Array_9_31_io_out_weight),
    .io_out_psum(PE_Array_9_31_io_out_psum)
  );
  basic_PE PE_Array_10_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_0_clock),
    .reset(PE_Array_10_0_reset),
    .io_in_activate(PE_Array_10_0_io_in_activate),
    .io_in_weight(PE_Array_10_0_io_in_weight),
    .io_in_psum(PE_Array_10_0_io_in_psum),
    .io_in_flow(PE_Array_10_0_io_in_flow),
    .io_in_shift(PE_Array_10_0_io_in_shift),
    .io_out_activate(PE_Array_10_0_io_out_activate),
    .io_out_weight(PE_Array_10_0_io_out_weight),
    .io_out_psum(PE_Array_10_0_io_out_psum)
  );
  basic_PE PE_Array_10_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_1_clock),
    .reset(PE_Array_10_1_reset),
    .io_in_activate(PE_Array_10_1_io_in_activate),
    .io_in_weight(PE_Array_10_1_io_in_weight),
    .io_in_psum(PE_Array_10_1_io_in_psum),
    .io_in_flow(PE_Array_10_1_io_in_flow),
    .io_in_shift(PE_Array_10_1_io_in_shift),
    .io_out_activate(PE_Array_10_1_io_out_activate),
    .io_out_weight(PE_Array_10_1_io_out_weight),
    .io_out_psum(PE_Array_10_1_io_out_psum)
  );
  basic_PE PE_Array_10_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_2_clock),
    .reset(PE_Array_10_2_reset),
    .io_in_activate(PE_Array_10_2_io_in_activate),
    .io_in_weight(PE_Array_10_2_io_in_weight),
    .io_in_psum(PE_Array_10_2_io_in_psum),
    .io_in_flow(PE_Array_10_2_io_in_flow),
    .io_in_shift(PE_Array_10_2_io_in_shift),
    .io_out_activate(PE_Array_10_2_io_out_activate),
    .io_out_weight(PE_Array_10_2_io_out_weight),
    .io_out_psum(PE_Array_10_2_io_out_psum)
  );
  basic_PE PE_Array_10_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_3_clock),
    .reset(PE_Array_10_3_reset),
    .io_in_activate(PE_Array_10_3_io_in_activate),
    .io_in_weight(PE_Array_10_3_io_in_weight),
    .io_in_psum(PE_Array_10_3_io_in_psum),
    .io_in_flow(PE_Array_10_3_io_in_flow),
    .io_in_shift(PE_Array_10_3_io_in_shift),
    .io_out_activate(PE_Array_10_3_io_out_activate),
    .io_out_weight(PE_Array_10_3_io_out_weight),
    .io_out_psum(PE_Array_10_3_io_out_psum)
  );
  basic_PE PE_Array_10_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_4_clock),
    .reset(PE_Array_10_4_reset),
    .io_in_activate(PE_Array_10_4_io_in_activate),
    .io_in_weight(PE_Array_10_4_io_in_weight),
    .io_in_psum(PE_Array_10_4_io_in_psum),
    .io_in_flow(PE_Array_10_4_io_in_flow),
    .io_in_shift(PE_Array_10_4_io_in_shift),
    .io_out_activate(PE_Array_10_4_io_out_activate),
    .io_out_weight(PE_Array_10_4_io_out_weight),
    .io_out_psum(PE_Array_10_4_io_out_psum)
  );
  basic_PE PE_Array_10_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_5_clock),
    .reset(PE_Array_10_5_reset),
    .io_in_activate(PE_Array_10_5_io_in_activate),
    .io_in_weight(PE_Array_10_5_io_in_weight),
    .io_in_psum(PE_Array_10_5_io_in_psum),
    .io_in_flow(PE_Array_10_5_io_in_flow),
    .io_in_shift(PE_Array_10_5_io_in_shift),
    .io_out_activate(PE_Array_10_5_io_out_activate),
    .io_out_weight(PE_Array_10_5_io_out_weight),
    .io_out_psum(PE_Array_10_5_io_out_psum)
  );
  basic_PE PE_Array_10_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_6_clock),
    .reset(PE_Array_10_6_reset),
    .io_in_activate(PE_Array_10_6_io_in_activate),
    .io_in_weight(PE_Array_10_6_io_in_weight),
    .io_in_psum(PE_Array_10_6_io_in_psum),
    .io_in_flow(PE_Array_10_6_io_in_flow),
    .io_in_shift(PE_Array_10_6_io_in_shift),
    .io_out_activate(PE_Array_10_6_io_out_activate),
    .io_out_weight(PE_Array_10_6_io_out_weight),
    .io_out_psum(PE_Array_10_6_io_out_psum)
  );
  basic_PE PE_Array_10_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_7_clock),
    .reset(PE_Array_10_7_reset),
    .io_in_activate(PE_Array_10_7_io_in_activate),
    .io_in_weight(PE_Array_10_7_io_in_weight),
    .io_in_psum(PE_Array_10_7_io_in_psum),
    .io_in_flow(PE_Array_10_7_io_in_flow),
    .io_in_shift(PE_Array_10_7_io_in_shift),
    .io_out_activate(PE_Array_10_7_io_out_activate),
    .io_out_weight(PE_Array_10_7_io_out_weight),
    .io_out_psum(PE_Array_10_7_io_out_psum)
  );
  basic_PE PE_Array_10_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_8_clock),
    .reset(PE_Array_10_8_reset),
    .io_in_activate(PE_Array_10_8_io_in_activate),
    .io_in_weight(PE_Array_10_8_io_in_weight),
    .io_in_psum(PE_Array_10_8_io_in_psum),
    .io_in_flow(PE_Array_10_8_io_in_flow),
    .io_in_shift(PE_Array_10_8_io_in_shift),
    .io_out_activate(PE_Array_10_8_io_out_activate),
    .io_out_weight(PE_Array_10_8_io_out_weight),
    .io_out_psum(PE_Array_10_8_io_out_psum)
  );
  basic_PE PE_Array_10_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_9_clock),
    .reset(PE_Array_10_9_reset),
    .io_in_activate(PE_Array_10_9_io_in_activate),
    .io_in_weight(PE_Array_10_9_io_in_weight),
    .io_in_psum(PE_Array_10_9_io_in_psum),
    .io_in_flow(PE_Array_10_9_io_in_flow),
    .io_in_shift(PE_Array_10_9_io_in_shift),
    .io_out_activate(PE_Array_10_9_io_out_activate),
    .io_out_weight(PE_Array_10_9_io_out_weight),
    .io_out_psum(PE_Array_10_9_io_out_psum)
  );
  basic_PE PE_Array_10_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_10_clock),
    .reset(PE_Array_10_10_reset),
    .io_in_activate(PE_Array_10_10_io_in_activate),
    .io_in_weight(PE_Array_10_10_io_in_weight),
    .io_in_psum(PE_Array_10_10_io_in_psum),
    .io_in_flow(PE_Array_10_10_io_in_flow),
    .io_in_shift(PE_Array_10_10_io_in_shift),
    .io_out_activate(PE_Array_10_10_io_out_activate),
    .io_out_weight(PE_Array_10_10_io_out_weight),
    .io_out_psum(PE_Array_10_10_io_out_psum)
  );
  basic_PE PE_Array_10_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_11_clock),
    .reset(PE_Array_10_11_reset),
    .io_in_activate(PE_Array_10_11_io_in_activate),
    .io_in_weight(PE_Array_10_11_io_in_weight),
    .io_in_psum(PE_Array_10_11_io_in_psum),
    .io_in_flow(PE_Array_10_11_io_in_flow),
    .io_in_shift(PE_Array_10_11_io_in_shift),
    .io_out_activate(PE_Array_10_11_io_out_activate),
    .io_out_weight(PE_Array_10_11_io_out_weight),
    .io_out_psum(PE_Array_10_11_io_out_psum)
  );
  basic_PE PE_Array_10_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_12_clock),
    .reset(PE_Array_10_12_reset),
    .io_in_activate(PE_Array_10_12_io_in_activate),
    .io_in_weight(PE_Array_10_12_io_in_weight),
    .io_in_psum(PE_Array_10_12_io_in_psum),
    .io_in_flow(PE_Array_10_12_io_in_flow),
    .io_in_shift(PE_Array_10_12_io_in_shift),
    .io_out_activate(PE_Array_10_12_io_out_activate),
    .io_out_weight(PE_Array_10_12_io_out_weight),
    .io_out_psum(PE_Array_10_12_io_out_psum)
  );
  basic_PE PE_Array_10_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_13_clock),
    .reset(PE_Array_10_13_reset),
    .io_in_activate(PE_Array_10_13_io_in_activate),
    .io_in_weight(PE_Array_10_13_io_in_weight),
    .io_in_psum(PE_Array_10_13_io_in_psum),
    .io_in_flow(PE_Array_10_13_io_in_flow),
    .io_in_shift(PE_Array_10_13_io_in_shift),
    .io_out_activate(PE_Array_10_13_io_out_activate),
    .io_out_weight(PE_Array_10_13_io_out_weight),
    .io_out_psum(PE_Array_10_13_io_out_psum)
  );
  basic_PE PE_Array_10_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_14_clock),
    .reset(PE_Array_10_14_reset),
    .io_in_activate(PE_Array_10_14_io_in_activate),
    .io_in_weight(PE_Array_10_14_io_in_weight),
    .io_in_psum(PE_Array_10_14_io_in_psum),
    .io_in_flow(PE_Array_10_14_io_in_flow),
    .io_in_shift(PE_Array_10_14_io_in_shift),
    .io_out_activate(PE_Array_10_14_io_out_activate),
    .io_out_weight(PE_Array_10_14_io_out_weight),
    .io_out_psum(PE_Array_10_14_io_out_psum)
  );
  basic_PE PE_Array_10_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_15_clock),
    .reset(PE_Array_10_15_reset),
    .io_in_activate(PE_Array_10_15_io_in_activate),
    .io_in_weight(PE_Array_10_15_io_in_weight),
    .io_in_psum(PE_Array_10_15_io_in_psum),
    .io_in_flow(PE_Array_10_15_io_in_flow),
    .io_in_shift(PE_Array_10_15_io_in_shift),
    .io_out_activate(PE_Array_10_15_io_out_activate),
    .io_out_weight(PE_Array_10_15_io_out_weight),
    .io_out_psum(PE_Array_10_15_io_out_psum)
  );
  basic_PE PE_Array_10_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_16_clock),
    .reset(PE_Array_10_16_reset),
    .io_in_activate(PE_Array_10_16_io_in_activate),
    .io_in_weight(PE_Array_10_16_io_in_weight),
    .io_in_psum(PE_Array_10_16_io_in_psum),
    .io_in_flow(PE_Array_10_16_io_in_flow),
    .io_in_shift(PE_Array_10_16_io_in_shift),
    .io_out_activate(PE_Array_10_16_io_out_activate),
    .io_out_weight(PE_Array_10_16_io_out_weight),
    .io_out_psum(PE_Array_10_16_io_out_psum)
  );
  basic_PE PE_Array_10_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_17_clock),
    .reset(PE_Array_10_17_reset),
    .io_in_activate(PE_Array_10_17_io_in_activate),
    .io_in_weight(PE_Array_10_17_io_in_weight),
    .io_in_psum(PE_Array_10_17_io_in_psum),
    .io_in_flow(PE_Array_10_17_io_in_flow),
    .io_in_shift(PE_Array_10_17_io_in_shift),
    .io_out_activate(PE_Array_10_17_io_out_activate),
    .io_out_weight(PE_Array_10_17_io_out_weight),
    .io_out_psum(PE_Array_10_17_io_out_psum)
  );
  basic_PE PE_Array_10_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_18_clock),
    .reset(PE_Array_10_18_reset),
    .io_in_activate(PE_Array_10_18_io_in_activate),
    .io_in_weight(PE_Array_10_18_io_in_weight),
    .io_in_psum(PE_Array_10_18_io_in_psum),
    .io_in_flow(PE_Array_10_18_io_in_flow),
    .io_in_shift(PE_Array_10_18_io_in_shift),
    .io_out_activate(PE_Array_10_18_io_out_activate),
    .io_out_weight(PE_Array_10_18_io_out_weight),
    .io_out_psum(PE_Array_10_18_io_out_psum)
  );
  basic_PE PE_Array_10_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_19_clock),
    .reset(PE_Array_10_19_reset),
    .io_in_activate(PE_Array_10_19_io_in_activate),
    .io_in_weight(PE_Array_10_19_io_in_weight),
    .io_in_psum(PE_Array_10_19_io_in_psum),
    .io_in_flow(PE_Array_10_19_io_in_flow),
    .io_in_shift(PE_Array_10_19_io_in_shift),
    .io_out_activate(PE_Array_10_19_io_out_activate),
    .io_out_weight(PE_Array_10_19_io_out_weight),
    .io_out_psum(PE_Array_10_19_io_out_psum)
  );
  basic_PE PE_Array_10_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_20_clock),
    .reset(PE_Array_10_20_reset),
    .io_in_activate(PE_Array_10_20_io_in_activate),
    .io_in_weight(PE_Array_10_20_io_in_weight),
    .io_in_psum(PE_Array_10_20_io_in_psum),
    .io_in_flow(PE_Array_10_20_io_in_flow),
    .io_in_shift(PE_Array_10_20_io_in_shift),
    .io_out_activate(PE_Array_10_20_io_out_activate),
    .io_out_weight(PE_Array_10_20_io_out_weight),
    .io_out_psum(PE_Array_10_20_io_out_psum)
  );
  basic_PE PE_Array_10_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_21_clock),
    .reset(PE_Array_10_21_reset),
    .io_in_activate(PE_Array_10_21_io_in_activate),
    .io_in_weight(PE_Array_10_21_io_in_weight),
    .io_in_psum(PE_Array_10_21_io_in_psum),
    .io_in_flow(PE_Array_10_21_io_in_flow),
    .io_in_shift(PE_Array_10_21_io_in_shift),
    .io_out_activate(PE_Array_10_21_io_out_activate),
    .io_out_weight(PE_Array_10_21_io_out_weight),
    .io_out_psum(PE_Array_10_21_io_out_psum)
  );
  basic_PE PE_Array_10_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_22_clock),
    .reset(PE_Array_10_22_reset),
    .io_in_activate(PE_Array_10_22_io_in_activate),
    .io_in_weight(PE_Array_10_22_io_in_weight),
    .io_in_psum(PE_Array_10_22_io_in_psum),
    .io_in_flow(PE_Array_10_22_io_in_flow),
    .io_in_shift(PE_Array_10_22_io_in_shift),
    .io_out_activate(PE_Array_10_22_io_out_activate),
    .io_out_weight(PE_Array_10_22_io_out_weight),
    .io_out_psum(PE_Array_10_22_io_out_psum)
  );
  basic_PE PE_Array_10_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_23_clock),
    .reset(PE_Array_10_23_reset),
    .io_in_activate(PE_Array_10_23_io_in_activate),
    .io_in_weight(PE_Array_10_23_io_in_weight),
    .io_in_psum(PE_Array_10_23_io_in_psum),
    .io_in_flow(PE_Array_10_23_io_in_flow),
    .io_in_shift(PE_Array_10_23_io_in_shift),
    .io_out_activate(PE_Array_10_23_io_out_activate),
    .io_out_weight(PE_Array_10_23_io_out_weight),
    .io_out_psum(PE_Array_10_23_io_out_psum)
  );
  basic_PE PE_Array_10_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_24_clock),
    .reset(PE_Array_10_24_reset),
    .io_in_activate(PE_Array_10_24_io_in_activate),
    .io_in_weight(PE_Array_10_24_io_in_weight),
    .io_in_psum(PE_Array_10_24_io_in_psum),
    .io_in_flow(PE_Array_10_24_io_in_flow),
    .io_in_shift(PE_Array_10_24_io_in_shift),
    .io_out_activate(PE_Array_10_24_io_out_activate),
    .io_out_weight(PE_Array_10_24_io_out_weight),
    .io_out_psum(PE_Array_10_24_io_out_psum)
  );
  basic_PE PE_Array_10_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_25_clock),
    .reset(PE_Array_10_25_reset),
    .io_in_activate(PE_Array_10_25_io_in_activate),
    .io_in_weight(PE_Array_10_25_io_in_weight),
    .io_in_psum(PE_Array_10_25_io_in_psum),
    .io_in_flow(PE_Array_10_25_io_in_flow),
    .io_in_shift(PE_Array_10_25_io_in_shift),
    .io_out_activate(PE_Array_10_25_io_out_activate),
    .io_out_weight(PE_Array_10_25_io_out_weight),
    .io_out_psum(PE_Array_10_25_io_out_psum)
  );
  basic_PE PE_Array_10_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_26_clock),
    .reset(PE_Array_10_26_reset),
    .io_in_activate(PE_Array_10_26_io_in_activate),
    .io_in_weight(PE_Array_10_26_io_in_weight),
    .io_in_psum(PE_Array_10_26_io_in_psum),
    .io_in_flow(PE_Array_10_26_io_in_flow),
    .io_in_shift(PE_Array_10_26_io_in_shift),
    .io_out_activate(PE_Array_10_26_io_out_activate),
    .io_out_weight(PE_Array_10_26_io_out_weight),
    .io_out_psum(PE_Array_10_26_io_out_psum)
  );
  basic_PE PE_Array_10_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_27_clock),
    .reset(PE_Array_10_27_reset),
    .io_in_activate(PE_Array_10_27_io_in_activate),
    .io_in_weight(PE_Array_10_27_io_in_weight),
    .io_in_psum(PE_Array_10_27_io_in_psum),
    .io_in_flow(PE_Array_10_27_io_in_flow),
    .io_in_shift(PE_Array_10_27_io_in_shift),
    .io_out_activate(PE_Array_10_27_io_out_activate),
    .io_out_weight(PE_Array_10_27_io_out_weight),
    .io_out_psum(PE_Array_10_27_io_out_psum)
  );
  basic_PE PE_Array_10_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_28_clock),
    .reset(PE_Array_10_28_reset),
    .io_in_activate(PE_Array_10_28_io_in_activate),
    .io_in_weight(PE_Array_10_28_io_in_weight),
    .io_in_psum(PE_Array_10_28_io_in_psum),
    .io_in_flow(PE_Array_10_28_io_in_flow),
    .io_in_shift(PE_Array_10_28_io_in_shift),
    .io_out_activate(PE_Array_10_28_io_out_activate),
    .io_out_weight(PE_Array_10_28_io_out_weight),
    .io_out_psum(PE_Array_10_28_io_out_psum)
  );
  basic_PE PE_Array_10_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_29_clock),
    .reset(PE_Array_10_29_reset),
    .io_in_activate(PE_Array_10_29_io_in_activate),
    .io_in_weight(PE_Array_10_29_io_in_weight),
    .io_in_psum(PE_Array_10_29_io_in_psum),
    .io_in_flow(PE_Array_10_29_io_in_flow),
    .io_in_shift(PE_Array_10_29_io_in_shift),
    .io_out_activate(PE_Array_10_29_io_out_activate),
    .io_out_weight(PE_Array_10_29_io_out_weight),
    .io_out_psum(PE_Array_10_29_io_out_psum)
  );
  basic_PE PE_Array_10_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_30_clock),
    .reset(PE_Array_10_30_reset),
    .io_in_activate(PE_Array_10_30_io_in_activate),
    .io_in_weight(PE_Array_10_30_io_in_weight),
    .io_in_psum(PE_Array_10_30_io_in_psum),
    .io_in_flow(PE_Array_10_30_io_in_flow),
    .io_in_shift(PE_Array_10_30_io_in_shift),
    .io_out_activate(PE_Array_10_30_io_out_activate),
    .io_out_weight(PE_Array_10_30_io_out_weight),
    .io_out_psum(PE_Array_10_30_io_out_psum)
  );
  basic_PE PE_Array_10_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_10_31_clock),
    .reset(PE_Array_10_31_reset),
    .io_in_activate(PE_Array_10_31_io_in_activate),
    .io_in_weight(PE_Array_10_31_io_in_weight),
    .io_in_psum(PE_Array_10_31_io_in_psum),
    .io_in_flow(PE_Array_10_31_io_in_flow),
    .io_in_shift(PE_Array_10_31_io_in_shift),
    .io_out_activate(PE_Array_10_31_io_out_activate),
    .io_out_weight(PE_Array_10_31_io_out_weight),
    .io_out_psum(PE_Array_10_31_io_out_psum)
  );
  basic_PE PE_Array_11_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_0_clock),
    .reset(PE_Array_11_0_reset),
    .io_in_activate(PE_Array_11_0_io_in_activate),
    .io_in_weight(PE_Array_11_0_io_in_weight),
    .io_in_psum(PE_Array_11_0_io_in_psum),
    .io_in_flow(PE_Array_11_0_io_in_flow),
    .io_in_shift(PE_Array_11_0_io_in_shift),
    .io_out_activate(PE_Array_11_0_io_out_activate),
    .io_out_weight(PE_Array_11_0_io_out_weight),
    .io_out_psum(PE_Array_11_0_io_out_psum)
  );
  basic_PE PE_Array_11_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_1_clock),
    .reset(PE_Array_11_1_reset),
    .io_in_activate(PE_Array_11_1_io_in_activate),
    .io_in_weight(PE_Array_11_1_io_in_weight),
    .io_in_psum(PE_Array_11_1_io_in_psum),
    .io_in_flow(PE_Array_11_1_io_in_flow),
    .io_in_shift(PE_Array_11_1_io_in_shift),
    .io_out_activate(PE_Array_11_1_io_out_activate),
    .io_out_weight(PE_Array_11_1_io_out_weight),
    .io_out_psum(PE_Array_11_1_io_out_psum)
  );
  basic_PE PE_Array_11_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_2_clock),
    .reset(PE_Array_11_2_reset),
    .io_in_activate(PE_Array_11_2_io_in_activate),
    .io_in_weight(PE_Array_11_2_io_in_weight),
    .io_in_psum(PE_Array_11_2_io_in_psum),
    .io_in_flow(PE_Array_11_2_io_in_flow),
    .io_in_shift(PE_Array_11_2_io_in_shift),
    .io_out_activate(PE_Array_11_2_io_out_activate),
    .io_out_weight(PE_Array_11_2_io_out_weight),
    .io_out_psum(PE_Array_11_2_io_out_psum)
  );
  basic_PE PE_Array_11_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_3_clock),
    .reset(PE_Array_11_3_reset),
    .io_in_activate(PE_Array_11_3_io_in_activate),
    .io_in_weight(PE_Array_11_3_io_in_weight),
    .io_in_psum(PE_Array_11_3_io_in_psum),
    .io_in_flow(PE_Array_11_3_io_in_flow),
    .io_in_shift(PE_Array_11_3_io_in_shift),
    .io_out_activate(PE_Array_11_3_io_out_activate),
    .io_out_weight(PE_Array_11_3_io_out_weight),
    .io_out_psum(PE_Array_11_3_io_out_psum)
  );
  basic_PE PE_Array_11_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_4_clock),
    .reset(PE_Array_11_4_reset),
    .io_in_activate(PE_Array_11_4_io_in_activate),
    .io_in_weight(PE_Array_11_4_io_in_weight),
    .io_in_psum(PE_Array_11_4_io_in_psum),
    .io_in_flow(PE_Array_11_4_io_in_flow),
    .io_in_shift(PE_Array_11_4_io_in_shift),
    .io_out_activate(PE_Array_11_4_io_out_activate),
    .io_out_weight(PE_Array_11_4_io_out_weight),
    .io_out_psum(PE_Array_11_4_io_out_psum)
  );
  basic_PE PE_Array_11_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_5_clock),
    .reset(PE_Array_11_5_reset),
    .io_in_activate(PE_Array_11_5_io_in_activate),
    .io_in_weight(PE_Array_11_5_io_in_weight),
    .io_in_psum(PE_Array_11_5_io_in_psum),
    .io_in_flow(PE_Array_11_5_io_in_flow),
    .io_in_shift(PE_Array_11_5_io_in_shift),
    .io_out_activate(PE_Array_11_5_io_out_activate),
    .io_out_weight(PE_Array_11_5_io_out_weight),
    .io_out_psum(PE_Array_11_5_io_out_psum)
  );
  basic_PE PE_Array_11_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_6_clock),
    .reset(PE_Array_11_6_reset),
    .io_in_activate(PE_Array_11_6_io_in_activate),
    .io_in_weight(PE_Array_11_6_io_in_weight),
    .io_in_psum(PE_Array_11_6_io_in_psum),
    .io_in_flow(PE_Array_11_6_io_in_flow),
    .io_in_shift(PE_Array_11_6_io_in_shift),
    .io_out_activate(PE_Array_11_6_io_out_activate),
    .io_out_weight(PE_Array_11_6_io_out_weight),
    .io_out_psum(PE_Array_11_6_io_out_psum)
  );
  basic_PE PE_Array_11_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_7_clock),
    .reset(PE_Array_11_7_reset),
    .io_in_activate(PE_Array_11_7_io_in_activate),
    .io_in_weight(PE_Array_11_7_io_in_weight),
    .io_in_psum(PE_Array_11_7_io_in_psum),
    .io_in_flow(PE_Array_11_7_io_in_flow),
    .io_in_shift(PE_Array_11_7_io_in_shift),
    .io_out_activate(PE_Array_11_7_io_out_activate),
    .io_out_weight(PE_Array_11_7_io_out_weight),
    .io_out_psum(PE_Array_11_7_io_out_psum)
  );
  basic_PE PE_Array_11_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_8_clock),
    .reset(PE_Array_11_8_reset),
    .io_in_activate(PE_Array_11_8_io_in_activate),
    .io_in_weight(PE_Array_11_8_io_in_weight),
    .io_in_psum(PE_Array_11_8_io_in_psum),
    .io_in_flow(PE_Array_11_8_io_in_flow),
    .io_in_shift(PE_Array_11_8_io_in_shift),
    .io_out_activate(PE_Array_11_8_io_out_activate),
    .io_out_weight(PE_Array_11_8_io_out_weight),
    .io_out_psum(PE_Array_11_8_io_out_psum)
  );
  basic_PE PE_Array_11_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_9_clock),
    .reset(PE_Array_11_9_reset),
    .io_in_activate(PE_Array_11_9_io_in_activate),
    .io_in_weight(PE_Array_11_9_io_in_weight),
    .io_in_psum(PE_Array_11_9_io_in_psum),
    .io_in_flow(PE_Array_11_9_io_in_flow),
    .io_in_shift(PE_Array_11_9_io_in_shift),
    .io_out_activate(PE_Array_11_9_io_out_activate),
    .io_out_weight(PE_Array_11_9_io_out_weight),
    .io_out_psum(PE_Array_11_9_io_out_psum)
  );
  basic_PE PE_Array_11_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_10_clock),
    .reset(PE_Array_11_10_reset),
    .io_in_activate(PE_Array_11_10_io_in_activate),
    .io_in_weight(PE_Array_11_10_io_in_weight),
    .io_in_psum(PE_Array_11_10_io_in_psum),
    .io_in_flow(PE_Array_11_10_io_in_flow),
    .io_in_shift(PE_Array_11_10_io_in_shift),
    .io_out_activate(PE_Array_11_10_io_out_activate),
    .io_out_weight(PE_Array_11_10_io_out_weight),
    .io_out_psum(PE_Array_11_10_io_out_psum)
  );
  basic_PE PE_Array_11_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_11_clock),
    .reset(PE_Array_11_11_reset),
    .io_in_activate(PE_Array_11_11_io_in_activate),
    .io_in_weight(PE_Array_11_11_io_in_weight),
    .io_in_psum(PE_Array_11_11_io_in_psum),
    .io_in_flow(PE_Array_11_11_io_in_flow),
    .io_in_shift(PE_Array_11_11_io_in_shift),
    .io_out_activate(PE_Array_11_11_io_out_activate),
    .io_out_weight(PE_Array_11_11_io_out_weight),
    .io_out_psum(PE_Array_11_11_io_out_psum)
  );
  basic_PE PE_Array_11_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_12_clock),
    .reset(PE_Array_11_12_reset),
    .io_in_activate(PE_Array_11_12_io_in_activate),
    .io_in_weight(PE_Array_11_12_io_in_weight),
    .io_in_psum(PE_Array_11_12_io_in_psum),
    .io_in_flow(PE_Array_11_12_io_in_flow),
    .io_in_shift(PE_Array_11_12_io_in_shift),
    .io_out_activate(PE_Array_11_12_io_out_activate),
    .io_out_weight(PE_Array_11_12_io_out_weight),
    .io_out_psum(PE_Array_11_12_io_out_psum)
  );
  basic_PE PE_Array_11_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_13_clock),
    .reset(PE_Array_11_13_reset),
    .io_in_activate(PE_Array_11_13_io_in_activate),
    .io_in_weight(PE_Array_11_13_io_in_weight),
    .io_in_psum(PE_Array_11_13_io_in_psum),
    .io_in_flow(PE_Array_11_13_io_in_flow),
    .io_in_shift(PE_Array_11_13_io_in_shift),
    .io_out_activate(PE_Array_11_13_io_out_activate),
    .io_out_weight(PE_Array_11_13_io_out_weight),
    .io_out_psum(PE_Array_11_13_io_out_psum)
  );
  basic_PE PE_Array_11_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_14_clock),
    .reset(PE_Array_11_14_reset),
    .io_in_activate(PE_Array_11_14_io_in_activate),
    .io_in_weight(PE_Array_11_14_io_in_weight),
    .io_in_psum(PE_Array_11_14_io_in_psum),
    .io_in_flow(PE_Array_11_14_io_in_flow),
    .io_in_shift(PE_Array_11_14_io_in_shift),
    .io_out_activate(PE_Array_11_14_io_out_activate),
    .io_out_weight(PE_Array_11_14_io_out_weight),
    .io_out_psum(PE_Array_11_14_io_out_psum)
  );
  basic_PE PE_Array_11_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_15_clock),
    .reset(PE_Array_11_15_reset),
    .io_in_activate(PE_Array_11_15_io_in_activate),
    .io_in_weight(PE_Array_11_15_io_in_weight),
    .io_in_psum(PE_Array_11_15_io_in_psum),
    .io_in_flow(PE_Array_11_15_io_in_flow),
    .io_in_shift(PE_Array_11_15_io_in_shift),
    .io_out_activate(PE_Array_11_15_io_out_activate),
    .io_out_weight(PE_Array_11_15_io_out_weight),
    .io_out_psum(PE_Array_11_15_io_out_psum)
  );
  basic_PE PE_Array_11_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_16_clock),
    .reset(PE_Array_11_16_reset),
    .io_in_activate(PE_Array_11_16_io_in_activate),
    .io_in_weight(PE_Array_11_16_io_in_weight),
    .io_in_psum(PE_Array_11_16_io_in_psum),
    .io_in_flow(PE_Array_11_16_io_in_flow),
    .io_in_shift(PE_Array_11_16_io_in_shift),
    .io_out_activate(PE_Array_11_16_io_out_activate),
    .io_out_weight(PE_Array_11_16_io_out_weight),
    .io_out_psum(PE_Array_11_16_io_out_psum)
  );
  basic_PE PE_Array_11_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_17_clock),
    .reset(PE_Array_11_17_reset),
    .io_in_activate(PE_Array_11_17_io_in_activate),
    .io_in_weight(PE_Array_11_17_io_in_weight),
    .io_in_psum(PE_Array_11_17_io_in_psum),
    .io_in_flow(PE_Array_11_17_io_in_flow),
    .io_in_shift(PE_Array_11_17_io_in_shift),
    .io_out_activate(PE_Array_11_17_io_out_activate),
    .io_out_weight(PE_Array_11_17_io_out_weight),
    .io_out_psum(PE_Array_11_17_io_out_psum)
  );
  basic_PE PE_Array_11_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_18_clock),
    .reset(PE_Array_11_18_reset),
    .io_in_activate(PE_Array_11_18_io_in_activate),
    .io_in_weight(PE_Array_11_18_io_in_weight),
    .io_in_psum(PE_Array_11_18_io_in_psum),
    .io_in_flow(PE_Array_11_18_io_in_flow),
    .io_in_shift(PE_Array_11_18_io_in_shift),
    .io_out_activate(PE_Array_11_18_io_out_activate),
    .io_out_weight(PE_Array_11_18_io_out_weight),
    .io_out_psum(PE_Array_11_18_io_out_psum)
  );
  basic_PE PE_Array_11_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_19_clock),
    .reset(PE_Array_11_19_reset),
    .io_in_activate(PE_Array_11_19_io_in_activate),
    .io_in_weight(PE_Array_11_19_io_in_weight),
    .io_in_psum(PE_Array_11_19_io_in_psum),
    .io_in_flow(PE_Array_11_19_io_in_flow),
    .io_in_shift(PE_Array_11_19_io_in_shift),
    .io_out_activate(PE_Array_11_19_io_out_activate),
    .io_out_weight(PE_Array_11_19_io_out_weight),
    .io_out_psum(PE_Array_11_19_io_out_psum)
  );
  basic_PE PE_Array_11_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_20_clock),
    .reset(PE_Array_11_20_reset),
    .io_in_activate(PE_Array_11_20_io_in_activate),
    .io_in_weight(PE_Array_11_20_io_in_weight),
    .io_in_psum(PE_Array_11_20_io_in_psum),
    .io_in_flow(PE_Array_11_20_io_in_flow),
    .io_in_shift(PE_Array_11_20_io_in_shift),
    .io_out_activate(PE_Array_11_20_io_out_activate),
    .io_out_weight(PE_Array_11_20_io_out_weight),
    .io_out_psum(PE_Array_11_20_io_out_psum)
  );
  basic_PE PE_Array_11_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_21_clock),
    .reset(PE_Array_11_21_reset),
    .io_in_activate(PE_Array_11_21_io_in_activate),
    .io_in_weight(PE_Array_11_21_io_in_weight),
    .io_in_psum(PE_Array_11_21_io_in_psum),
    .io_in_flow(PE_Array_11_21_io_in_flow),
    .io_in_shift(PE_Array_11_21_io_in_shift),
    .io_out_activate(PE_Array_11_21_io_out_activate),
    .io_out_weight(PE_Array_11_21_io_out_weight),
    .io_out_psum(PE_Array_11_21_io_out_psum)
  );
  basic_PE PE_Array_11_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_22_clock),
    .reset(PE_Array_11_22_reset),
    .io_in_activate(PE_Array_11_22_io_in_activate),
    .io_in_weight(PE_Array_11_22_io_in_weight),
    .io_in_psum(PE_Array_11_22_io_in_psum),
    .io_in_flow(PE_Array_11_22_io_in_flow),
    .io_in_shift(PE_Array_11_22_io_in_shift),
    .io_out_activate(PE_Array_11_22_io_out_activate),
    .io_out_weight(PE_Array_11_22_io_out_weight),
    .io_out_psum(PE_Array_11_22_io_out_psum)
  );
  basic_PE PE_Array_11_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_23_clock),
    .reset(PE_Array_11_23_reset),
    .io_in_activate(PE_Array_11_23_io_in_activate),
    .io_in_weight(PE_Array_11_23_io_in_weight),
    .io_in_psum(PE_Array_11_23_io_in_psum),
    .io_in_flow(PE_Array_11_23_io_in_flow),
    .io_in_shift(PE_Array_11_23_io_in_shift),
    .io_out_activate(PE_Array_11_23_io_out_activate),
    .io_out_weight(PE_Array_11_23_io_out_weight),
    .io_out_psum(PE_Array_11_23_io_out_psum)
  );
  basic_PE PE_Array_11_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_24_clock),
    .reset(PE_Array_11_24_reset),
    .io_in_activate(PE_Array_11_24_io_in_activate),
    .io_in_weight(PE_Array_11_24_io_in_weight),
    .io_in_psum(PE_Array_11_24_io_in_psum),
    .io_in_flow(PE_Array_11_24_io_in_flow),
    .io_in_shift(PE_Array_11_24_io_in_shift),
    .io_out_activate(PE_Array_11_24_io_out_activate),
    .io_out_weight(PE_Array_11_24_io_out_weight),
    .io_out_psum(PE_Array_11_24_io_out_psum)
  );
  basic_PE PE_Array_11_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_25_clock),
    .reset(PE_Array_11_25_reset),
    .io_in_activate(PE_Array_11_25_io_in_activate),
    .io_in_weight(PE_Array_11_25_io_in_weight),
    .io_in_psum(PE_Array_11_25_io_in_psum),
    .io_in_flow(PE_Array_11_25_io_in_flow),
    .io_in_shift(PE_Array_11_25_io_in_shift),
    .io_out_activate(PE_Array_11_25_io_out_activate),
    .io_out_weight(PE_Array_11_25_io_out_weight),
    .io_out_psum(PE_Array_11_25_io_out_psum)
  );
  basic_PE PE_Array_11_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_26_clock),
    .reset(PE_Array_11_26_reset),
    .io_in_activate(PE_Array_11_26_io_in_activate),
    .io_in_weight(PE_Array_11_26_io_in_weight),
    .io_in_psum(PE_Array_11_26_io_in_psum),
    .io_in_flow(PE_Array_11_26_io_in_flow),
    .io_in_shift(PE_Array_11_26_io_in_shift),
    .io_out_activate(PE_Array_11_26_io_out_activate),
    .io_out_weight(PE_Array_11_26_io_out_weight),
    .io_out_psum(PE_Array_11_26_io_out_psum)
  );
  basic_PE PE_Array_11_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_27_clock),
    .reset(PE_Array_11_27_reset),
    .io_in_activate(PE_Array_11_27_io_in_activate),
    .io_in_weight(PE_Array_11_27_io_in_weight),
    .io_in_psum(PE_Array_11_27_io_in_psum),
    .io_in_flow(PE_Array_11_27_io_in_flow),
    .io_in_shift(PE_Array_11_27_io_in_shift),
    .io_out_activate(PE_Array_11_27_io_out_activate),
    .io_out_weight(PE_Array_11_27_io_out_weight),
    .io_out_psum(PE_Array_11_27_io_out_psum)
  );
  basic_PE PE_Array_11_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_28_clock),
    .reset(PE_Array_11_28_reset),
    .io_in_activate(PE_Array_11_28_io_in_activate),
    .io_in_weight(PE_Array_11_28_io_in_weight),
    .io_in_psum(PE_Array_11_28_io_in_psum),
    .io_in_flow(PE_Array_11_28_io_in_flow),
    .io_in_shift(PE_Array_11_28_io_in_shift),
    .io_out_activate(PE_Array_11_28_io_out_activate),
    .io_out_weight(PE_Array_11_28_io_out_weight),
    .io_out_psum(PE_Array_11_28_io_out_psum)
  );
  basic_PE PE_Array_11_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_29_clock),
    .reset(PE_Array_11_29_reset),
    .io_in_activate(PE_Array_11_29_io_in_activate),
    .io_in_weight(PE_Array_11_29_io_in_weight),
    .io_in_psum(PE_Array_11_29_io_in_psum),
    .io_in_flow(PE_Array_11_29_io_in_flow),
    .io_in_shift(PE_Array_11_29_io_in_shift),
    .io_out_activate(PE_Array_11_29_io_out_activate),
    .io_out_weight(PE_Array_11_29_io_out_weight),
    .io_out_psum(PE_Array_11_29_io_out_psum)
  );
  basic_PE PE_Array_11_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_30_clock),
    .reset(PE_Array_11_30_reset),
    .io_in_activate(PE_Array_11_30_io_in_activate),
    .io_in_weight(PE_Array_11_30_io_in_weight),
    .io_in_psum(PE_Array_11_30_io_in_psum),
    .io_in_flow(PE_Array_11_30_io_in_flow),
    .io_in_shift(PE_Array_11_30_io_in_shift),
    .io_out_activate(PE_Array_11_30_io_out_activate),
    .io_out_weight(PE_Array_11_30_io_out_weight),
    .io_out_psum(PE_Array_11_30_io_out_psum)
  );
  basic_PE PE_Array_11_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_11_31_clock),
    .reset(PE_Array_11_31_reset),
    .io_in_activate(PE_Array_11_31_io_in_activate),
    .io_in_weight(PE_Array_11_31_io_in_weight),
    .io_in_psum(PE_Array_11_31_io_in_psum),
    .io_in_flow(PE_Array_11_31_io_in_flow),
    .io_in_shift(PE_Array_11_31_io_in_shift),
    .io_out_activate(PE_Array_11_31_io_out_activate),
    .io_out_weight(PE_Array_11_31_io_out_weight),
    .io_out_psum(PE_Array_11_31_io_out_psum)
  );
  basic_PE PE_Array_12_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_0_clock),
    .reset(PE_Array_12_0_reset),
    .io_in_activate(PE_Array_12_0_io_in_activate),
    .io_in_weight(PE_Array_12_0_io_in_weight),
    .io_in_psum(PE_Array_12_0_io_in_psum),
    .io_in_flow(PE_Array_12_0_io_in_flow),
    .io_in_shift(PE_Array_12_0_io_in_shift),
    .io_out_activate(PE_Array_12_0_io_out_activate),
    .io_out_weight(PE_Array_12_0_io_out_weight),
    .io_out_psum(PE_Array_12_0_io_out_psum)
  );
  basic_PE PE_Array_12_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_1_clock),
    .reset(PE_Array_12_1_reset),
    .io_in_activate(PE_Array_12_1_io_in_activate),
    .io_in_weight(PE_Array_12_1_io_in_weight),
    .io_in_psum(PE_Array_12_1_io_in_psum),
    .io_in_flow(PE_Array_12_1_io_in_flow),
    .io_in_shift(PE_Array_12_1_io_in_shift),
    .io_out_activate(PE_Array_12_1_io_out_activate),
    .io_out_weight(PE_Array_12_1_io_out_weight),
    .io_out_psum(PE_Array_12_1_io_out_psum)
  );
  basic_PE PE_Array_12_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_2_clock),
    .reset(PE_Array_12_2_reset),
    .io_in_activate(PE_Array_12_2_io_in_activate),
    .io_in_weight(PE_Array_12_2_io_in_weight),
    .io_in_psum(PE_Array_12_2_io_in_psum),
    .io_in_flow(PE_Array_12_2_io_in_flow),
    .io_in_shift(PE_Array_12_2_io_in_shift),
    .io_out_activate(PE_Array_12_2_io_out_activate),
    .io_out_weight(PE_Array_12_2_io_out_weight),
    .io_out_psum(PE_Array_12_2_io_out_psum)
  );
  basic_PE PE_Array_12_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_3_clock),
    .reset(PE_Array_12_3_reset),
    .io_in_activate(PE_Array_12_3_io_in_activate),
    .io_in_weight(PE_Array_12_3_io_in_weight),
    .io_in_psum(PE_Array_12_3_io_in_psum),
    .io_in_flow(PE_Array_12_3_io_in_flow),
    .io_in_shift(PE_Array_12_3_io_in_shift),
    .io_out_activate(PE_Array_12_3_io_out_activate),
    .io_out_weight(PE_Array_12_3_io_out_weight),
    .io_out_psum(PE_Array_12_3_io_out_psum)
  );
  basic_PE PE_Array_12_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_4_clock),
    .reset(PE_Array_12_4_reset),
    .io_in_activate(PE_Array_12_4_io_in_activate),
    .io_in_weight(PE_Array_12_4_io_in_weight),
    .io_in_psum(PE_Array_12_4_io_in_psum),
    .io_in_flow(PE_Array_12_4_io_in_flow),
    .io_in_shift(PE_Array_12_4_io_in_shift),
    .io_out_activate(PE_Array_12_4_io_out_activate),
    .io_out_weight(PE_Array_12_4_io_out_weight),
    .io_out_psum(PE_Array_12_4_io_out_psum)
  );
  basic_PE PE_Array_12_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_5_clock),
    .reset(PE_Array_12_5_reset),
    .io_in_activate(PE_Array_12_5_io_in_activate),
    .io_in_weight(PE_Array_12_5_io_in_weight),
    .io_in_psum(PE_Array_12_5_io_in_psum),
    .io_in_flow(PE_Array_12_5_io_in_flow),
    .io_in_shift(PE_Array_12_5_io_in_shift),
    .io_out_activate(PE_Array_12_5_io_out_activate),
    .io_out_weight(PE_Array_12_5_io_out_weight),
    .io_out_psum(PE_Array_12_5_io_out_psum)
  );
  basic_PE PE_Array_12_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_6_clock),
    .reset(PE_Array_12_6_reset),
    .io_in_activate(PE_Array_12_6_io_in_activate),
    .io_in_weight(PE_Array_12_6_io_in_weight),
    .io_in_psum(PE_Array_12_6_io_in_psum),
    .io_in_flow(PE_Array_12_6_io_in_flow),
    .io_in_shift(PE_Array_12_6_io_in_shift),
    .io_out_activate(PE_Array_12_6_io_out_activate),
    .io_out_weight(PE_Array_12_6_io_out_weight),
    .io_out_psum(PE_Array_12_6_io_out_psum)
  );
  basic_PE PE_Array_12_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_7_clock),
    .reset(PE_Array_12_7_reset),
    .io_in_activate(PE_Array_12_7_io_in_activate),
    .io_in_weight(PE_Array_12_7_io_in_weight),
    .io_in_psum(PE_Array_12_7_io_in_psum),
    .io_in_flow(PE_Array_12_7_io_in_flow),
    .io_in_shift(PE_Array_12_7_io_in_shift),
    .io_out_activate(PE_Array_12_7_io_out_activate),
    .io_out_weight(PE_Array_12_7_io_out_weight),
    .io_out_psum(PE_Array_12_7_io_out_psum)
  );
  basic_PE PE_Array_12_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_8_clock),
    .reset(PE_Array_12_8_reset),
    .io_in_activate(PE_Array_12_8_io_in_activate),
    .io_in_weight(PE_Array_12_8_io_in_weight),
    .io_in_psum(PE_Array_12_8_io_in_psum),
    .io_in_flow(PE_Array_12_8_io_in_flow),
    .io_in_shift(PE_Array_12_8_io_in_shift),
    .io_out_activate(PE_Array_12_8_io_out_activate),
    .io_out_weight(PE_Array_12_8_io_out_weight),
    .io_out_psum(PE_Array_12_8_io_out_psum)
  );
  basic_PE PE_Array_12_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_9_clock),
    .reset(PE_Array_12_9_reset),
    .io_in_activate(PE_Array_12_9_io_in_activate),
    .io_in_weight(PE_Array_12_9_io_in_weight),
    .io_in_psum(PE_Array_12_9_io_in_psum),
    .io_in_flow(PE_Array_12_9_io_in_flow),
    .io_in_shift(PE_Array_12_9_io_in_shift),
    .io_out_activate(PE_Array_12_9_io_out_activate),
    .io_out_weight(PE_Array_12_9_io_out_weight),
    .io_out_psum(PE_Array_12_9_io_out_psum)
  );
  basic_PE PE_Array_12_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_10_clock),
    .reset(PE_Array_12_10_reset),
    .io_in_activate(PE_Array_12_10_io_in_activate),
    .io_in_weight(PE_Array_12_10_io_in_weight),
    .io_in_psum(PE_Array_12_10_io_in_psum),
    .io_in_flow(PE_Array_12_10_io_in_flow),
    .io_in_shift(PE_Array_12_10_io_in_shift),
    .io_out_activate(PE_Array_12_10_io_out_activate),
    .io_out_weight(PE_Array_12_10_io_out_weight),
    .io_out_psum(PE_Array_12_10_io_out_psum)
  );
  basic_PE PE_Array_12_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_11_clock),
    .reset(PE_Array_12_11_reset),
    .io_in_activate(PE_Array_12_11_io_in_activate),
    .io_in_weight(PE_Array_12_11_io_in_weight),
    .io_in_psum(PE_Array_12_11_io_in_psum),
    .io_in_flow(PE_Array_12_11_io_in_flow),
    .io_in_shift(PE_Array_12_11_io_in_shift),
    .io_out_activate(PE_Array_12_11_io_out_activate),
    .io_out_weight(PE_Array_12_11_io_out_weight),
    .io_out_psum(PE_Array_12_11_io_out_psum)
  );
  basic_PE PE_Array_12_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_12_clock),
    .reset(PE_Array_12_12_reset),
    .io_in_activate(PE_Array_12_12_io_in_activate),
    .io_in_weight(PE_Array_12_12_io_in_weight),
    .io_in_psum(PE_Array_12_12_io_in_psum),
    .io_in_flow(PE_Array_12_12_io_in_flow),
    .io_in_shift(PE_Array_12_12_io_in_shift),
    .io_out_activate(PE_Array_12_12_io_out_activate),
    .io_out_weight(PE_Array_12_12_io_out_weight),
    .io_out_psum(PE_Array_12_12_io_out_psum)
  );
  basic_PE PE_Array_12_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_13_clock),
    .reset(PE_Array_12_13_reset),
    .io_in_activate(PE_Array_12_13_io_in_activate),
    .io_in_weight(PE_Array_12_13_io_in_weight),
    .io_in_psum(PE_Array_12_13_io_in_psum),
    .io_in_flow(PE_Array_12_13_io_in_flow),
    .io_in_shift(PE_Array_12_13_io_in_shift),
    .io_out_activate(PE_Array_12_13_io_out_activate),
    .io_out_weight(PE_Array_12_13_io_out_weight),
    .io_out_psum(PE_Array_12_13_io_out_psum)
  );
  basic_PE PE_Array_12_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_14_clock),
    .reset(PE_Array_12_14_reset),
    .io_in_activate(PE_Array_12_14_io_in_activate),
    .io_in_weight(PE_Array_12_14_io_in_weight),
    .io_in_psum(PE_Array_12_14_io_in_psum),
    .io_in_flow(PE_Array_12_14_io_in_flow),
    .io_in_shift(PE_Array_12_14_io_in_shift),
    .io_out_activate(PE_Array_12_14_io_out_activate),
    .io_out_weight(PE_Array_12_14_io_out_weight),
    .io_out_psum(PE_Array_12_14_io_out_psum)
  );
  basic_PE PE_Array_12_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_15_clock),
    .reset(PE_Array_12_15_reset),
    .io_in_activate(PE_Array_12_15_io_in_activate),
    .io_in_weight(PE_Array_12_15_io_in_weight),
    .io_in_psum(PE_Array_12_15_io_in_psum),
    .io_in_flow(PE_Array_12_15_io_in_flow),
    .io_in_shift(PE_Array_12_15_io_in_shift),
    .io_out_activate(PE_Array_12_15_io_out_activate),
    .io_out_weight(PE_Array_12_15_io_out_weight),
    .io_out_psum(PE_Array_12_15_io_out_psum)
  );
  basic_PE PE_Array_12_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_16_clock),
    .reset(PE_Array_12_16_reset),
    .io_in_activate(PE_Array_12_16_io_in_activate),
    .io_in_weight(PE_Array_12_16_io_in_weight),
    .io_in_psum(PE_Array_12_16_io_in_psum),
    .io_in_flow(PE_Array_12_16_io_in_flow),
    .io_in_shift(PE_Array_12_16_io_in_shift),
    .io_out_activate(PE_Array_12_16_io_out_activate),
    .io_out_weight(PE_Array_12_16_io_out_weight),
    .io_out_psum(PE_Array_12_16_io_out_psum)
  );
  basic_PE PE_Array_12_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_17_clock),
    .reset(PE_Array_12_17_reset),
    .io_in_activate(PE_Array_12_17_io_in_activate),
    .io_in_weight(PE_Array_12_17_io_in_weight),
    .io_in_psum(PE_Array_12_17_io_in_psum),
    .io_in_flow(PE_Array_12_17_io_in_flow),
    .io_in_shift(PE_Array_12_17_io_in_shift),
    .io_out_activate(PE_Array_12_17_io_out_activate),
    .io_out_weight(PE_Array_12_17_io_out_weight),
    .io_out_psum(PE_Array_12_17_io_out_psum)
  );
  basic_PE PE_Array_12_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_18_clock),
    .reset(PE_Array_12_18_reset),
    .io_in_activate(PE_Array_12_18_io_in_activate),
    .io_in_weight(PE_Array_12_18_io_in_weight),
    .io_in_psum(PE_Array_12_18_io_in_psum),
    .io_in_flow(PE_Array_12_18_io_in_flow),
    .io_in_shift(PE_Array_12_18_io_in_shift),
    .io_out_activate(PE_Array_12_18_io_out_activate),
    .io_out_weight(PE_Array_12_18_io_out_weight),
    .io_out_psum(PE_Array_12_18_io_out_psum)
  );
  basic_PE PE_Array_12_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_19_clock),
    .reset(PE_Array_12_19_reset),
    .io_in_activate(PE_Array_12_19_io_in_activate),
    .io_in_weight(PE_Array_12_19_io_in_weight),
    .io_in_psum(PE_Array_12_19_io_in_psum),
    .io_in_flow(PE_Array_12_19_io_in_flow),
    .io_in_shift(PE_Array_12_19_io_in_shift),
    .io_out_activate(PE_Array_12_19_io_out_activate),
    .io_out_weight(PE_Array_12_19_io_out_weight),
    .io_out_psum(PE_Array_12_19_io_out_psum)
  );
  basic_PE PE_Array_12_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_20_clock),
    .reset(PE_Array_12_20_reset),
    .io_in_activate(PE_Array_12_20_io_in_activate),
    .io_in_weight(PE_Array_12_20_io_in_weight),
    .io_in_psum(PE_Array_12_20_io_in_psum),
    .io_in_flow(PE_Array_12_20_io_in_flow),
    .io_in_shift(PE_Array_12_20_io_in_shift),
    .io_out_activate(PE_Array_12_20_io_out_activate),
    .io_out_weight(PE_Array_12_20_io_out_weight),
    .io_out_psum(PE_Array_12_20_io_out_psum)
  );
  basic_PE PE_Array_12_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_21_clock),
    .reset(PE_Array_12_21_reset),
    .io_in_activate(PE_Array_12_21_io_in_activate),
    .io_in_weight(PE_Array_12_21_io_in_weight),
    .io_in_psum(PE_Array_12_21_io_in_psum),
    .io_in_flow(PE_Array_12_21_io_in_flow),
    .io_in_shift(PE_Array_12_21_io_in_shift),
    .io_out_activate(PE_Array_12_21_io_out_activate),
    .io_out_weight(PE_Array_12_21_io_out_weight),
    .io_out_psum(PE_Array_12_21_io_out_psum)
  );
  basic_PE PE_Array_12_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_22_clock),
    .reset(PE_Array_12_22_reset),
    .io_in_activate(PE_Array_12_22_io_in_activate),
    .io_in_weight(PE_Array_12_22_io_in_weight),
    .io_in_psum(PE_Array_12_22_io_in_psum),
    .io_in_flow(PE_Array_12_22_io_in_flow),
    .io_in_shift(PE_Array_12_22_io_in_shift),
    .io_out_activate(PE_Array_12_22_io_out_activate),
    .io_out_weight(PE_Array_12_22_io_out_weight),
    .io_out_psum(PE_Array_12_22_io_out_psum)
  );
  basic_PE PE_Array_12_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_23_clock),
    .reset(PE_Array_12_23_reset),
    .io_in_activate(PE_Array_12_23_io_in_activate),
    .io_in_weight(PE_Array_12_23_io_in_weight),
    .io_in_psum(PE_Array_12_23_io_in_psum),
    .io_in_flow(PE_Array_12_23_io_in_flow),
    .io_in_shift(PE_Array_12_23_io_in_shift),
    .io_out_activate(PE_Array_12_23_io_out_activate),
    .io_out_weight(PE_Array_12_23_io_out_weight),
    .io_out_psum(PE_Array_12_23_io_out_psum)
  );
  basic_PE PE_Array_12_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_24_clock),
    .reset(PE_Array_12_24_reset),
    .io_in_activate(PE_Array_12_24_io_in_activate),
    .io_in_weight(PE_Array_12_24_io_in_weight),
    .io_in_psum(PE_Array_12_24_io_in_psum),
    .io_in_flow(PE_Array_12_24_io_in_flow),
    .io_in_shift(PE_Array_12_24_io_in_shift),
    .io_out_activate(PE_Array_12_24_io_out_activate),
    .io_out_weight(PE_Array_12_24_io_out_weight),
    .io_out_psum(PE_Array_12_24_io_out_psum)
  );
  basic_PE PE_Array_12_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_25_clock),
    .reset(PE_Array_12_25_reset),
    .io_in_activate(PE_Array_12_25_io_in_activate),
    .io_in_weight(PE_Array_12_25_io_in_weight),
    .io_in_psum(PE_Array_12_25_io_in_psum),
    .io_in_flow(PE_Array_12_25_io_in_flow),
    .io_in_shift(PE_Array_12_25_io_in_shift),
    .io_out_activate(PE_Array_12_25_io_out_activate),
    .io_out_weight(PE_Array_12_25_io_out_weight),
    .io_out_psum(PE_Array_12_25_io_out_psum)
  );
  basic_PE PE_Array_12_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_26_clock),
    .reset(PE_Array_12_26_reset),
    .io_in_activate(PE_Array_12_26_io_in_activate),
    .io_in_weight(PE_Array_12_26_io_in_weight),
    .io_in_psum(PE_Array_12_26_io_in_psum),
    .io_in_flow(PE_Array_12_26_io_in_flow),
    .io_in_shift(PE_Array_12_26_io_in_shift),
    .io_out_activate(PE_Array_12_26_io_out_activate),
    .io_out_weight(PE_Array_12_26_io_out_weight),
    .io_out_psum(PE_Array_12_26_io_out_psum)
  );
  basic_PE PE_Array_12_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_27_clock),
    .reset(PE_Array_12_27_reset),
    .io_in_activate(PE_Array_12_27_io_in_activate),
    .io_in_weight(PE_Array_12_27_io_in_weight),
    .io_in_psum(PE_Array_12_27_io_in_psum),
    .io_in_flow(PE_Array_12_27_io_in_flow),
    .io_in_shift(PE_Array_12_27_io_in_shift),
    .io_out_activate(PE_Array_12_27_io_out_activate),
    .io_out_weight(PE_Array_12_27_io_out_weight),
    .io_out_psum(PE_Array_12_27_io_out_psum)
  );
  basic_PE PE_Array_12_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_28_clock),
    .reset(PE_Array_12_28_reset),
    .io_in_activate(PE_Array_12_28_io_in_activate),
    .io_in_weight(PE_Array_12_28_io_in_weight),
    .io_in_psum(PE_Array_12_28_io_in_psum),
    .io_in_flow(PE_Array_12_28_io_in_flow),
    .io_in_shift(PE_Array_12_28_io_in_shift),
    .io_out_activate(PE_Array_12_28_io_out_activate),
    .io_out_weight(PE_Array_12_28_io_out_weight),
    .io_out_psum(PE_Array_12_28_io_out_psum)
  );
  basic_PE PE_Array_12_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_29_clock),
    .reset(PE_Array_12_29_reset),
    .io_in_activate(PE_Array_12_29_io_in_activate),
    .io_in_weight(PE_Array_12_29_io_in_weight),
    .io_in_psum(PE_Array_12_29_io_in_psum),
    .io_in_flow(PE_Array_12_29_io_in_flow),
    .io_in_shift(PE_Array_12_29_io_in_shift),
    .io_out_activate(PE_Array_12_29_io_out_activate),
    .io_out_weight(PE_Array_12_29_io_out_weight),
    .io_out_psum(PE_Array_12_29_io_out_psum)
  );
  basic_PE PE_Array_12_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_30_clock),
    .reset(PE_Array_12_30_reset),
    .io_in_activate(PE_Array_12_30_io_in_activate),
    .io_in_weight(PE_Array_12_30_io_in_weight),
    .io_in_psum(PE_Array_12_30_io_in_psum),
    .io_in_flow(PE_Array_12_30_io_in_flow),
    .io_in_shift(PE_Array_12_30_io_in_shift),
    .io_out_activate(PE_Array_12_30_io_out_activate),
    .io_out_weight(PE_Array_12_30_io_out_weight),
    .io_out_psum(PE_Array_12_30_io_out_psum)
  );
  basic_PE PE_Array_12_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_12_31_clock),
    .reset(PE_Array_12_31_reset),
    .io_in_activate(PE_Array_12_31_io_in_activate),
    .io_in_weight(PE_Array_12_31_io_in_weight),
    .io_in_psum(PE_Array_12_31_io_in_psum),
    .io_in_flow(PE_Array_12_31_io_in_flow),
    .io_in_shift(PE_Array_12_31_io_in_shift),
    .io_out_activate(PE_Array_12_31_io_out_activate),
    .io_out_weight(PE_Array_12_31_io_out_weight),
    .io_out_psum(PE_Array_12_31_io_out_psum)
  );
  basic_PE PE_Array_13_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_0_clock),
    .reset(PE_Array_13_0_reset),
    .io_in_activate(PE_Array_13_0_io_in_activate),
    .io_in_weight(PE_Array_13_0_io_in_weight),
    .io_in_psum(PE_Array_13_0_io_in_psum),
    .io_in_flow(PE_Array_13_0_io_in_flow),
    .io_in_shift(PE_Array_13_0_io_in_shift),
    .io_out_activate(PE_Array_13_0_io_out_activate),
    .io_out_weight(PE_Array_13_0_io_out_weight),
    .io_out_psum(PE_Array_13_0_io_out_psum)
  );
  basic_PE PE_Array_13_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_1_clock),
    .reset(PE_Array_13_1_reset),
    .io_in_activate(PE_Array_13_1_io_in_activate),
    .io_in_weight(PE_Array_13_1_io_in_weight),
    .io_in_psum(PE_Array_13_1_io_in_psum),
    .io_in_flow(PE_Array_13_1_io_in_flow),
    .io_in_shift(PE_Array_13_1_io_in_shift),
    .io_out_activate(PE_Array_13_1_io_out_activate),
    .io_out_weight(PE_Array_13_1_io_out_weight),
    .io_out_psum(PE_Array_13_1_io_out_psum)
  );
  basic_PE PE_Array_13_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_2_clock),
    .reset(PE_Array_13_2_reset),
    .io_in_activate(PE_Array_13_2_io_in_activate),
    .io_in_weight(PE_Array_13_2_io_in_weight),
    .io_in_psum(PE_Array_13_2_io_in_psum),
    .io_in_flow(PE_Array_13_2_io_in_flow),
    .io_in_shift(PE_Array_13_2_io_in_shift),
    .io_out_activate(PE_Array_13_2_io_out_activate),
    .io_out_weight(PE_Array_13_2_io_out_weight),
    .io_out_psum(PE_Array_13_2_io_out_psum)
  );
  basic_PE PE_Array_13_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_3_clock),
    .reset(PE_Array_13_3_reset),
    .io_in_activate(PE_Array_13_3_io_in_activate),
    .io_in_weight(PE_Array_13_3_io_in_weight),
    .io_in_psum(PE_Array_13_3_io_in_psum),
    .io_in_flow(PE_Array_13_3_io_in_flow),
    .io_in_shift(PE_Array_13_3_io_in_shift),
    .io_out_activate(PE_Array_13_3_io_out_activate),
    .io_out_weight(PE_Array_13_3_io_out_weight),
    .io_out_psum(PE_Array_13_3_io_out_psum)
  );
  basic_PE PE_Array_13_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_4_clock),
    .reset(PE_Array_13_4_reset),
    .io_in_activate(PE_Array_13_4_io_in_activate),
    .io_in_weight(PE_Array_13_4_io_in_weight),
    .io_in_psum(PE_Array_13_4_io_in_psum),
    .io_in_flow(PE_Array_13_4_io_in_flow),
    .io_in_shift(PE_Array_13_4_io_in_shift),
    .io_out_activate(PE_Array_13_4_io_out_activate),
    .io_out_weight(PE_Array_13_4_io_out_weight),
    .io_out_psum(PE_Array_13_4_io_out_psum)
  );
  basic_PE PE_Array_13_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_5_clock),
    .reset(PE_Array_13_5_reset),
    .io_in_activate(PE_Array_13_5_io_in_activate),
    .io_in_weight(PE_Array_13_5_io_in_weight),
    .io_in_psum(PE_Array_13_5_io_in_psum),
    .io_in_flow(PE_Array_13_5_io_in_flow),
    .io_in_shift(PE_Array_13_5_io_in_shift),
    .io_out_activate(PE_Array_13_5_io_out_activate),
    .io_out_weight(PE_Array_13_5_io_out_weight),
    .io_out_psum(PE_Array_13_5_io_out_psum)
  );
  basic_PE PE_Array_13_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_6_clock),
    .reset(PE_Array_13_6_reset),
    .io_in_activate(PE_Array_13_6_io_in_activate),
    .io_in_weight(PE_Array_13_6_io_in_weight),
    .io_in_psum(PE_Array_13_6_io_in_psum),
    .io_in_flow(PE_Array_13_6_io_in_flow),
    .io_in_shift(PE_Array_13_6_io_in_shift),
    .io_out_activate(PE_Array_13_6_io_out_activate),
    .io_out_weight(PE_Array_13_6_io_out_weight),
    .io_out_psum(PE_Array_13_6_io_out_psum)
  );
  basic_PE PE_Array_13_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_7_clock),
    .reset(PE_Array_13_7_reset),
    .io_in_activate(PE_Array_13_7_io_in_activate),
    .io_in_weight(PE_Array_13_7_io_in_weight),
    .io_in_psum(PE_Array_13_7_io_in_psum),
    .io_in_flow(PE_Array_13_7_io_in_flow),
    .io_in_shift(PE_Array_13_7_io_in_shift),
    .io_out_activate(PE_Array_13_7_io_out_activate),
    .io_out_weight(PE_Array_13_7_io_out_weight),
    .io_out_psum(PE_Array_13_7_io_out_psum)
  );
  basic_PE PE_Array_13_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_8_clock),
    .reset(PE_Array_13_8_reset),
    .io_in_activate(PE_Array_13_8_io_in_activate),
    .io_in_weight(PE_Array_13_8_io_in_weight),
    .io_in_psum(PE_Array_13_8_io_in_psum),
    .io_in_flow(PE_Array_13_8_io_in_flow),
    .io_in_shift(PE_Array_13_8_io_in_shift),
    .io_out_activate(PE_Array_13_8_io_out_activate),
    .io_out_weight(PE_Array_13_8_io_out_weight),
    .io_out_psum(PE_Array_13_8_io_out_psum)
  );
  basic_PE PE_Array_13_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_9_clock),
    .reset(PE_Array_13_9_reset),
    .io_in_activate(PE_Array_13_9_io_in_activate),
    .io_in_weight(PE_Array_13_9_io_in_weight),
    .io_in_psum(PE_Array_13_9_io_in_psum),
    .io_in_flow(PE_Array_13_9_io_in_flow),
    .io_in_shift(PE_Array_13_9_io_in_shift),
    .io_out_activate(PE_Array_13_9_io_out_activate),
    .io_out_weight(PE_Array_13_9_io_out_weight),
    .io_out_psum(PE_Array_13_9_io_out_psum)
  );
  basic_PE PE_Array_13_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_10_clock),
    .reset(PE_Array_13_10_reset),
    .io_in_activate(PE_Array_13_10_io_in_activate),
    .io_in_weight(PE_Array_13_10_io_in_weight),
    .io_in_psum(PE_Array_13_10_io_in_psum),
    .io_in_flow(PE_Array_13_10_io_in_flow),
    .io_in_shift(PE_Array_13_10_io_in_shift),
    .io_out_activate(PE_Array_13_10_io_out_activate),
    .io_out_weight(PE_Array_13_10_io_out_weight),
    .io_out_psum(PE_Array_13_10_io_out_psum)
  );
  basic_PE PE_Array_13_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_11_clock),
    .reset(PE_Array_13_11_reset),
    .io_in_activate(PE_Array_13_11_io_in_activate),
    .io_in_weight(PE_Array_13_11_io_in_weight),
    .io_in_psum(PE_Array_13_11_io_in_psum),
    .io_in_flow(PE_Array_13_11_io_in_flow),
    .io_in_shift(PE_Array_13_11_io_in_shift),
    .io_out_activate(PE_Array_13_11_io_out_activate),
    .io_out_weight(PE_Array_13_11_io_out_weight),
    .io_out_psum(PE_Array_13_11_io_out_psum)
  );
  basic_PE PE_Array_13_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_12_clock),
    .reset(PE_Array_13_12_reset),
    .io_in_activate(PE_Array_13_12_io_in_activate),
    .io_in_weight(PE_Array_13_12_io_in_weight),
    .io_in_psum(PE_Array_13_12_io_in_psum),
    .io_in_flow(PE_Array_13_12_io_in_flow),
    .io_in_shift(PE_Array_13_12_io_in_shift),
    .io_out_activate(PE_Array_13_12_io_out_activate),
    .io_out_weight(PE_Array_13_12_io_out_weight),
    .io_out_psum(PE_Array_13_12_io_out_psum)
  );
  basic_PE PE_Array_13_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_13_clock),
    .reset(PE_Array_13_13_reset),
    .io_in_activate(PE_Array_13_13_io_in_activate),
    .io_in_weight(PE_Array_13_13_io_in_weight),
    .io_in_psum(PE_Array_13_13_io_in_psum),
    .io_in_flow(PE_Array_13_13_io_in_flow),
    .io_in_shift(PE_Array_13_13_io_in_shift),
    .io_out_activate(PE_Array_13_13_io_out_activate),
    .io_out_weight(PE_Array_13_13_io_out_weight),
    .io_out_psum(PE_Array_13_13_io_out_psum)
  );
  basic_PE PE_Array_13_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_14_clock),
    .reset(PE_Array_13_14_reset),
    .io_in_activate(PE_Array_13_14_io_in_activate),
    .io_in_weight(PE_Array_13_14_io_in_weight),
    .io_in_psum(PE_Array_13_14_io_in_psum),
    .io_in_flow(PE_Array_13_14_io_in_flow),
    .io_in_shift(PE_Array_13_14_io_in_shift),
    .io_out_activate(PE_Array_13_14_io_out_activate),
    .io_out_weight(PE_Array_13_14_io_out_weight),
    .io_out_psum(PE_Array_13_14_io_out_psum)
  );
  basic_PE PE_Array_13_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_15_clock),
    .reset(PE_Array_13_15_reset),
    .io_in_activate(PE_Array_13_15_io_in_activate),
    .io_in_weight(PE_Array_13_15_io_in_weight),
    .io_in_psum(PE_Array_13_15_io_in_psum),
    .io_in_flow(PE_Array_13_15_io_in_flow),
    .io_in_shift(PE_Array_13_15_io_in_shift),
    .io_out_activate(PE_Array_13_15_io_out_activate),
    .io_out_weight(PE_Array_13_15_io_out_weight),
    .io_out_psum(PE_Array_13_15_io_out_psum)
  );
  basic_PE PE_Array_13_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_16_clock),
    .reset(PE_Array_13_16_reset),
    .io_in_activate(PE_Array_13_16_io_in_activate),
    .io_in_weight(PE_Array_13_16_io_in_weight),
    .io_in_psum(PE_Array_13_16_io_in_psum),
    .io_in_flow(PE_Array_13_16_io_in_flow),
    .io_in_shift(PE_Array_13_16_io_in_shift),
    .io_out_activate(PE_Array_13_16_io_out_activate),
    .io_out_weight(PE_Array_13_16_io_out_weight),
    .io_out_psum(PE_Array_13_16_io_out_psum)
  );
  basic_PE PE_Array_13_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_17_clock),
    .reset(PE_Array_13_17_reset),
    .io_in_activate(PE_Array_13_17_io_in_activate),
    .io_in_weight(PE_Array_13_17_io_in_weight),
    .io_in_psum(PE_Array_13_17_io_in_psum),
    .io_in_flow(PE_Array_13_17_io_in_flow),
    .io_in_shift(PE_Array_13_17_io_in_shift),
    .io_out_activate(PE_Array_13_17_io_out_activate),
    .io_out_weight(PE_Array_13_17_io_out_weight),
    .io_out_psum(PE_Array_13_17_io_out_psum)
  );
  basic_PE PE_Array_13_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_18_clock),
    .reset(PE_Array_13_18_reset),
    .io_in_activate(PE_Array_13_18_io_in_activate),
    .io_in_weight(PE_Array_13_18_io_in_weight),
    .io_in_psum(PE_Array_13_18_io_in_psum),
    .io_in_flow(PE_Array_13_18_io_in_flow),
    .io_in_shift(PE_Array_13_18_io_in_shift),
    .io_out_activate(PE_Array_13_18_io_out_activate),
    .io_out_weight(PE_Array_13_18_io_out_weight),
    .io_out_psum(PE_Array_13_18_io_out_psum)
  );
  basic_PE PE_Array_13_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_19_clock),
    .reset(PE_Array_13_19_reset),
    .io_in_activate(PE_Array_13_19_io_in_activate),
    .io_in_weight(PE_Array_13_19_io_in_weight),
    .io_in_psum(PE_Array_13_19_io_in_psum),
    .io_in_flow(PE_Array_13_19_io_in_flow),
    .io_in_shift(PE_Array_13_19_io_in_shift),
    .io_out_activate(PE_Array_13_19_io_out_activate),
    .io_out_weight(PE_Array_13_19_io_out_weight),
    .io_out_psum(PE_Array_13_19_io_out_psum)
  );
  basic_PE PE_Array_13_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_20_clock),
    .reset(PE_Array_13_20_reset),
    .io_in_activate(PE_Array_13_20_io_in_activate),
    .io_in_weight(PE_Array_13_20_io_in_weight),
    .io_in_psum(PE_Array_13_20_io_in_psum),
    .io_in_flow(PE_Array_13_20_io_in_flow),
    .io_in_shift(PE_Array_13_20_io_in_shift),
    .io_out_activate(PE_Array_13_20_io_out_activate),
    .io_out_weight(PE_Array_13_20_io_out_weight),
    .io_out_psum(PE_Array_13_20_io_out_psum)
  );
  basic_PE PE_Array_13_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_21_clock),
    .reset(PE_Array_13_21_reset),
    .io_in_activate(PE_Array_13_21_io_in_activate),
    .io_in_weight(PE_Array_13_21_io_in_weight),
    .io_in_psum(PE_Array_13_21_io_in_psum),
    .io_in_flow(PE_Array_13_21_io_in_flow),
    .io_in_shift(PE_Array_13_21_io_in_shift),
    .io_out_activate(PE_Array_13_21_io_out_activate),
    .io_out_weight(PE_Array_13_21_io_out_weight),
    .io_out_psum(PE_Array_13_21_io_out_psum)
  );
  basic_PE PE_Array_13_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_22_clock),
    .reset(PE_Array_13_22_reset),
    .io_in_activate(PE_Array_13_22_io_in_activate),
    .io_in_weight(PE_Array_13_22_io_in_weight),
    .io_in_psum(PE_Array_13_22_io_in_psum),
    .io_in_flow(PE_Array_13_22_io_in_flow),
    .io_in_shift(PE_Array_13_22_io_in_shift),
    .io_out_activate(PE_Array_13_22_io_out_activate),
    .io_out_weight(PE_Array_13_22_io_out_weight),
    .io_out_psum(PE_Array_13_22_io_out_psum)
  );
  basic_PE PE_Array_13_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_23_clock),
    .reset(PE_Array_13_23_reset),
    .io_in_activate(PE_Array_13_23_io_in_activate),
    .io_in_weight(PE_Array_13_23_io_in_weight),
    .io_in_psum(PE_Array_13_23_io_in_psum),
    .io_in_flow(PE_Array_13_23_io_in_flow),
    .io_in_shift(PE_Array_13_23_io_in_shift),
    .io_out_activate(PE_Array_13_23_io_out_activate),
    .io_out_weight(PE_Array_13_23_io_out_weight),
    .io_out_psum(PE_Array_13_23_io_out_psum)
  );
  basic_PE PE_Array_13_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_24_clock),
    .reset(PE_Array_13_24_reset),
    .io_in_activate(PE_Array_13_24_io_in_activate),
    .io_in_weight(PE_Array_13_24_io_in_weight),
    .io_in_psum(PE_Array_13_24_io_in_psum),
    .io_in_flow(PE_Array_13_24_io_in_flow),
    .io_in_shift(PE_Array_13_24_io_in_shift),
    .io_out_activate(PE_Array_13_24_io_out_activate),
    .io_out_weight(PE_Array_13_24_io_out_weight),
    .io_out_psum(PE_Array_13_24_io_out_psum)
  );
  basic_PE PE_Array_13_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_25_clock),
    .reset(PE_Array_13_25_reset),
    .io_in_activate(PE_Array_13_25_io_in_activate),
    .io_in_weight(PE_Array_13_25_io_in_weight),
    .io_in_psum(PE_Array_13_25_io_in_psum),
    .io_in_flow(PE_Array_13_25_io_in_flow),
    .io_in_shift(PE_Array_13_25_io_in_shift),
    .io_out_activate(PE_Array_13_25_io_out_activate),
    .io_out_weight(PE_Array_13_25_io_out_weight),
    .io_out_psum(PE_Array_13_25_io_out_psum)
  );
  basic_PE PE_Array_13_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_26_clock),
    .reset(PE_Array_13_26_reset),
    .io_in_activate(PE_Array_13_26_io_in_activate),
    .io_in_weight(PE_Array_13_26_io_in_weight),
    .io_in_psum(PE_Array_13_26_io_in_psum),
    .io_in_flow(PE_Array_13_26_io_in_flow),
    .io_in_shift(PE_Array_13_26_io_in_shift),
    .io_out_activate(PE_Array_13_26_io_out_activate),
    .io_out_weight(PE_Array_13_26_io_out_weight),
    .io_out_psum(PE_Array_13_26_io_out_psum)
  );
  basic_PE PE_Array_13_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_27_clock),
    .reset(PE_Array_13_27_reset),
    .io_in_activate(PE_Array_13_27_io_in_activate),
    .io_in_weight(PE_Array_13_27_io_in_weight),
    .io_in_psum(PE_Array_13_27_io_in_psum),
    .io_in_flow(PE_Array_13_27_io_in_flow),
    .io_in_shift(PE_Array_13_27_io_in_shift),
    .io_out_activate(PE_Array_13_27_io_out_activate),
    .io_out_weight(PE_Array_13_27_io_out_weight),
    .io_out_psum(PE_Array_13_27_io_out_psum)
  );
  basic_PE PE_Array_13_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_28_clock),
    .reset(PE_Array_13_28_reset),
    .io_in_activate(PE_Array_13_28_io_in_activate),
    .io_in_weight(PE_Array_13_28_io_in_weight),
    .io_in_psum(PE_Array_13_28_io_in_psum),
    .io_in_flow(PE_Array_13_28_io_in_flow),
    .io_in_shift(PE_Array_13_28_io_in_shift),
    .io_out_activate(PE_Array_13_28_io_out_activate),
    .io_out_weight(PE_Array_13_28_io_out_weight),
    .io_out_psum(PE_Array_13_28_io_out_psum)
  );
  basic_PE PE_Array_13_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_29_clock),
    .reset(PE_Array_13_29_reset),
    .io_in_activate(PE_Array_13_29_io_in_activate),
    .io_in_weight(PE_Array_13_29_io_in_weight),
    .io_in_psum(PE_Array_13_29_io_in_psum),
    .io_in_flow(PE_Array_13_29_io_in_flow),
    .io_in_shift(PE_Array_13_29_io_in_shift),
    .io_out_activate(PE_Array_13_29_io_out_activate),
    .io_out_weight(PE_Array_13_29_io_out_weight),
    .io_out_psum(PE_Array_13_29_io_out_psum)
  );
  basic_PE PE_Array_13_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_30_clock),
    .reset(PE_Array_13_30_reset),
    .io_in_activate(PE_Array_13_30_io_in_activate),
    .io_in_weight(PE_Array_13_30_io_in_weight),
    .io_in_psum(PE_Array_13_30_io_in_psum),
    .io_in_flow(PE_Array_13_30_io_in_flow),
    .io_in_shift(PE_Array_13_30_io_in_shift),
    .io_out_activate(PE_Array_13_30_io_out_activate),
    .io_out_weight(PE_Array_13_30_io_out_weight),
    .io_out_psum(PE_Array_13_30_io_out_psum)
  );
  basic_PE PE_Array_13_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_13_31_clock),
    .reset(PE_Array_13_31_reset),
    .io_in_activate(PE_Array_13_31_io_in_activate),
    .io_in_weight(PE_Array_13_31_io_in_weight),
    .io_in_psum(PE_Array_13_31_io_in_psum),
    .io_in_flow(PE_Array_13_31_io_in_flow),
    .io_in_shift(PE_Array_13_31_io_in_shift),
    .io_out_activate(PE_Array_13_31_io_out_activate),
    .io_out_weight(PE_Array_13_31_io_out_weight),
    .io_out_psum(PE_Array_13_31_io_out_psum)
  );
  basic_PE PE_Array_14_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_0_clock),
    .reset(PE_Array_14_0_reset),
    .io_in_activate(PE_Array_14_0_io_in_activate),
    .io_in_weight(PE_Array_14_0_io_in_weight),
    .io_in_psum(PE_Array_14_0_io_in_psum),
    .io_in_flow(PE_Array_14_0_io_in_flow),
    .io_in_shift(PE_Array_14_0_io_in_shift),
    .io_out_activate(PE_Array_14_0_io_out_activate),
    .io_out_weight(PE_Array_14_0_io_out_weight),
    .io_out_psum(PE_Array_14_0_io_out_psum)
  );
  basic_PE PE_Array_14_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_1_clock),
    .reset(PE_Array_14_1_reset),
    .io_in_activate(PE_Array_14_1_io_in_activate),
    .io_in_weight(PE_Array_14_1_io_in_weight),
    .io_in_psum(PE_Array_14_1_io_in_psum),
    .io_in_flow(PE_Array_14_1_io_in_flow),
    .io_in_shift(PE_Array_14_1_io_in_shift),
    .io_out_activate(PE_Array_14_1_io_out_activate),
    .io_out_weight(PE_Array_14_1_io_out_weight),
    .io_out_psum(PE_Array_14_1_io_out_psum)
  );
  basic_PE PE_Array_14_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_2_clock),
    .reset(PE_Array_14_2_reset),
    .io_in_activate(PE_Array_14_2_io_in_activate),
    .io_in_weight(PE_Array_14_2_io_in_weight),
    .io_in_psum(PE_Array_14_2_io_in_psum),
    .io_in_flow(PE_Array_14_2_io_in_flow),
    .io_in_shift(PE_Array_14_2_io_in_shift),
    .io_out_activate(PE_Array_14_2_io_out_activate),
    .io_out_weight(PE_Array_14_2_io_out_weight),
    .io_out_psum(PE_Array_14_2_io_out_psum)
  );
  basic_PE PE_Array_14_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_3_clock),
    .reset(PE_Array_14_3_reset),
    .io_in_activate(PE_Array_14_3_io_in_activate),
    .io_in_weight(PE_Array_14_3_io_in_weight),
    .io_in_psum(PE_Array_14_3_io_in_psum),
    .io_in_flow(PE_Array_14_3_io_in_flow),
    .io_in_shift(PE_Array_14_3_io_in_shift),
    .io_out_activate(PE_Array_14_3_io_out_activate),
    .io_out_weight(PE_Array_14_3_io_out_weight),
    .io_out_psum(PE_Array_14_3_io_out_psum)
  );
  basic_PE PE_Array_14_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_4_clock),
    .reset(PE_Array_14_4_reset),
    .io_in_activate(PE_Array_14_4_io_in_activate),
    .io_in_weight(PE_Array_14_4_io_in_weight),
    .io_in_psum(PE_Array_14_4_io_in_psum),
    .io_in_flow(PE_Array_14_4_io_in_flow),
    .io_in_shift(PE_Array_14_4_io_in_shift),
    .io_out_activate(PE_Array_14_4_io_out_activate),
    .io_out_weight(PE_Array_14_4_io_out_weight),
    .io_out_psum(PE_Array_14_4_io_out_psum)
  );
  basic_PE PE_Array_14_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_5_clock),
    .reset(PE_Array_14_5_reset),
    .io_in_activate(PE_Array_14_5_io_in_activate),
    .io_in_weight(PE_Array_14_5_io_in_weight),
    .io_in_psum(PE_Array_14_5_io_in_psum),
    .io_in_flow(PE_Array_14_5_io_in_flow),
    .io_in_shift(PE_Array_14_5_io_in_shift),
    .io_out_activate(PE_Array_14_5_io_out_activate),
    .io_out_weight(PE_Array_14_5_io_out_weight),
    .io_out_psum(PE_Array_14_5_io_out_psum)
  );
  basic_PE PE_Array_14_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_6_clock),
    .reset(PE_Array_14_6_reset),
    .io_in_activate(PE_Array_14_6_io_in_activate),
    .io_in_weight(PE_Array_14_6_io_in_weight),
    .io_in_psum(PE_Array_14_6_io_in_psum),
    .io_in_flow(PE_Array_14_6_io_in_flow),
    .io_in_shift(PE_Array_14_6_io_in_shift),
    .io_out_activate(PE_Array_14_6_io_out_activate),
    .io_out_weight(PE_Array_14_6_io_out_weight),
    .io_out_psum(PE_Array_14_6_io_out_psum)
  );
  basic_PE PE_Array_14_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_7_clock),
    .reset(PE_Array_14_7_reset),
    .io_in_activate(PE_Array_14_7_io_in_activate),
    .io_in_weight(PE_Array_14_7_io_in_weight),
    .io_in_psum(PE_Array_14_7_io_in_psum),
    .io_in_flow(PE_Array_14_7_io_in_flow),
    .io_in_shift(PE_Array_14_7_io_in_shift),
    .io_out_activate(PE_Array_14_7_io_out_activate),
    .io_out_weight(PE_Array_14_7_io_out_weight),
    .io_out_psum(PE_Array_14_7_io_out_psum)
  );
  basic_PE PE_Array_14_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_8_clock),
    .reset(PE_Array_14_8_reset),
    .io_in_activate(PE_Array_14_8_io_in_activate),
    .io_in_weight(PE_Array_14_8_io_in_weight),
    .io_in_psum(PE_Array_14_8_io_in_psum),
    .io_in_flow(PE_Array_14_8_io_in_flow),
    .io_in_shift(PE_Array_14_8_io_in_shift),
    .io_out_activate(PE_Array_14_8_io_out_activate),
    .io_out_weight(PE_Array_14_8_io_out_weight),
    .io_out_psum(PE_Array_14_8_io_out_psum)
  );
  basic_PE PE_Array_14_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_9_clock),
    .reset(PE_Array_14_9_reset),
    .io_in_activate(PE_Array_14_9_io_in_activate),
    .io_in_weight(PE_Array_14_9_io_in_weight),
    .io_in_psum(PE_Array_14_9_io_in_psum),
    .io_in_flow(PE_Array_14_9_io_in_flow),
    .io_in_shift(PE_Array_14_9_io_in_shift),
    .io_out_activate(PE_Array_14_9_io_out_activate),
    .io_out_weight(PE_Array_14_9_io_out_weight),
    .io_out_psum(PE_Array_14_9_io_out_psum)
  );
  basic_PE PE_Array_14_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_10_clock),
    .reset(PE_Array_14_10_reset),
    .io_in_activate(PE_Array_14_10_io_in_activate),
    .io_in_weight(PE_Array_14_10_io_in_weight),
    .io_in_psum(PE_Array_14_10_io_in_psum),
    .io_in_flow(PE_Array_14_10_io_in_flow),
    .io_in_shift(PE_Array_14_10_io_in_shift),
    .io_out_activate(PE_Array_14_10_io_out_activate),
    .io_out_weight(PE_Array_14_10_io_out_weight),
    .io_out_psum(PE_Array_14_10_io_out_psum)
  );
  basic_PE PE_Array_14_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_11_clock),
    .reset(PE_Array_14_11_reset),
    .io_in_activate(PE_Array_14_11_io_in_activate),
    .io_in_weight(PE_Array_14_11_io_in_weight),
    .io_in_psum(PE_Array_14_11_io_in_psum),
    .io_in_flow(PE_Array_14_11_io_in_flow),
    .io_in_shift(PE_Array_14_11_io_in_shift),
    .io_out_activate(PE_Array_14_11_io_out_activate),
    .io_out_weight(PE_Array_14_11_io_out_weight),
    .io_out_psum(PE_Array_14_11_io_out_psum)
  );
  basic_PE PE_Array_14_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_12_clock),
    .reset(PE_Array_14_12_reset),
    .io_in_activate(PE_Array_14_12_io_in_activate),
    .io_in_weight(PE_Array_14_12_io_in_weight),
    .io_in_psum(PE_Array_14_12_io_in_psum),
    .io_in_flow(PE_Array_14_12_io_in_flow),
    .io_in_shift(PE_Array_14_12_io_in_shift),
    .io_out_activate(PE_Array_14_12_io_out_activate),
    .io_out_weight(PE_Array_14_12_io_out_weight),
    .io_out_psum(PE_Array_14_12_io_out_psum)
  );
  basic_PE PE_Array_14_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_13_clock),
    .reset(PE_Array_14_13_reset),
    .io_in_activate(PE_Array_14_13_io_in_activate),
    .io_in_weight(PE_Array_14_13_io_in_weight),
    .io_in_psum(PE_Array_14_13_io_in_psum),
    .io_in_flow(PE_Array_14_13_io_in_flow),
    .io_in_shift(PE_Array_14_13_io_in_shift),
    .io_out_activate(PE_Array_14_13_io_out_activate),
    .io_out_weight(PE_Array_14_13_io_out_weight),
    .io_out_psum(PE_Array_14_13_io_out_psum)
  );
  basic_PE PE_Array_14_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_14_clock),
    .reset(PE_Array_14_14_reset),
    .io_in_activate(PE_Array_14_14_io_in_activate),
    .io_in_weight(PE_Array_14_14_io_in_weight),
    .io_in_psum(PE_Array_14_14_io_in_psum),
    .io_in_flow(PE_Array_14_14_io_in_flow),
    .io_in_shift(PE_Array_14_14_io_in_shift),
    .io_out_activate(PE_Array_14_14_io_out_activate),
    .io_out_weight(PE_Array_14_14_io_out_weight),
    .io_out_psum(PE_Array_14_14_io_out_psum)
  );
  basic_PE PE_Array_14_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_15_clock),
    .reset(PE_Array_14_15_reset),
    .io_in_activate(PE_Array_14_15_io_in_activate),
    .io_in_weight(PE_Array_14_15_io_in_weight),
    .io_in_psum(PE_Array_14_15_io_in_psum),
    .io_in_flow(PE_Array_14_15_io_in_flow),
    .io_in_shift(PE_Array_14_15_io_in_shift),
    .io_out_activate(PE_Array_14_15_io_out_activate),
    .io_out_weight(PE_Array_14_15_io_out_weight),
    .io_out_psum(PE_Array_14_15_io_out_psum)
  );
  basic_PE PE_Array_14_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_16_clock),
    .reset(PE_Array_14_16_reset),
    .io_in_activate(PE_Array_14_16_io_in_activate),
    .io_in_weight(PE_Array_14_16_io_in_weight),
    .io_in_psum(PE_Array_14_16_io_in_psum),
    .io_in_flow(PE_Array_14_16_io_in_flow),
    .io_in_shift(PE_Array_14_16_io_in_shift),
    .io_out_activate(PE_Array_14_16_io_out_activate),
    .io_out_weight(PE_Array_14_16_io_out_weight),
    .io_out_psum(PE_Array_14_16_io_out_psum)
  );
  basic_PE PE_Array_14_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_17_clock),
    .reset(PE_Array_14_17_reset),
    .io_in_activate(PE_Array_14_17_io_in_activate),
    .io_in_weight(PE_Array_14_17_io_in_weight),
    .io_in_psum(PE_Array_14_17_io_in_psum),
    .io_in_flow(PE_Array_14_17_io_in_flow),
    .io_in_shift(PE_Array_14_17_io_in_shift),
    .io_out_activate(PE_Array_14_17_io_out_activate),
    .io_out_weight(PE_Array_14_17_io_out_weight),
    .io_out_psum(PE_Array_14_17_io_out_psum)
  );
  basic_PE PE_Array_14_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_18_clock),
    .reset(PE_Array_14_18_reset),
    .io_in_activate(PE_Array_14_18_io_in_activate),
    .io_in_weight(PE_Array_14_18_io_in_weight),
    .io_in_psum(PE_Array_14_18_io_in_psum),
    .io_in_flow(PE_Array_14_18_io_in_flow),
    .io_in_shift(PE_Array_14_18_io_in_shift),
    .io_out_activate(PE_Array_14_18_io_out_activate),
    .io_out_weight(PE_Array_14_18_io_out_weight),
    .io_out_psum(PE_Array_14_18_io_out_psum)
  );
  basic_PE PE_Array_14_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_19_clock),
    .reset(PE_Array_14_19_reset),
    .io_in_activate(PE_Array_14_19_io_in_activate),
    .io_in_weight(PE_Array_14_19_io_in_weight),
    .io_in_psum(PE_Array_14_19_io_in_psum),
    .io_in_flow(PE_Array_14_19_io_in_flow),
    .io_in_shift(PE_Array_14_19_io_in_shift),
    .io_out_activate(PE_Array_14_19_io_out_activate),
    .io_out_weight(PE_Array_14_19_io_out_weight),
    .io_out_psum(PE_Array_14_19_io_out_psum)
  );
  basic_PE PE_Array_14_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_20_clock),
    .reset(PE_Array_14_20_reset),
    .io_in_activate(PE_Array_14_20_io_in_activate),
    .io_in_weight(PE_Array_14_20_io_in_weight),
    .io_in_psum(PE_Array_14_20_io_in_psum),
    .io_in_flow(PE_Array_14_20_io_in_flow),
    .io_in_shift(PE_Array_14_20_io_in_shift),
    .io_out_activate(PE_Array_14_20_io_out_activate),
    .io_out_weight(PE_Array_14_20_io_out_weight),
    .io_out_psum(PE_Array_14_20_io_out_psum)
  );
  basic_PE PE_Array_14_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_21_clock),
    .reset(PE_Array_14_21_reset),
    .io_in_activate(PE_Array_14_21_io_in_activate),
    .io_in_weight(PE_Array_14_21_io_in_weight),
    .io_in_psum(PE_Array_14_21_io_in_psum),
    .io_in_flow(PE_Array_14_21_io_in_flow),
    .io_in_shift(PE_Array_14_21_io_in_shift),
    .io_out_activate(PE_Array_14_21_io_out_activate),
    .io_out_weight(PE_Array_14_21_io_out_weight),
    .io_out_psum(PE_Array_14_21_io_out_psum)
  );
  basic_PE PE_Array_14_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_22_clock),
    .reset(PE_Array_14_22_reset),
    .io_in_activate(PE_Array_14_22_io_in_activate),
    .io_in_weight(PE_Array_14_22_io_in_weight),
    .io_in_psum(PE_Array_14_22_io_in_psum),
    .io_in_flow(PE_Array_14_22_io_in_flow),
    .io_in_shift(PE_Array_14_22_io_in_shift),
    .io_out_activate(PE_Array_14_22_io_out_activate),
    .io_out_weight(PE_Array_14_22_io_out_weight),
    .io_out_psum(PE_Array_14_22_io_out_psum)
  );
  basic_PE PE_Array_14_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_23_clock),
    .reset(PE_Array_14_23_reset),
    .io_in_activate(PE_Array_14_23_io_in_activate),
    .io_in_weight(PE_Array_14_23_io_in_weight),
    .io_in_psum(PE_Array_14_23_io_in_psum),
    .io_in_flow(PE_Array_14_23_io_in_flow),
    .io_in_shift(PE_Array_14_23_io_in_shift),
    .io_out_activate(PE_Array_14_23_io_out_activate),
    .io_out_weight(PE_Array_14_23_io_out_weight),
    .io_out_psum(PE_Array_14_23_io_out_psum)
  );
  basic_PE PE_Array_14_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_24_clock),
    .reset(PE_Array_14_24_reset),
    .io_in_activate(PE_Array_14_24_io_in_activate),
    .io_in_weight(PE_Array_14_24_io_in_weight),
    .io_in_psum(PE_Array_14_24_io_in_psum),
    .io_in_flow(PE_Array_14_24_io_in_flow),
    .io_in_shift(PE_Array_14_24_io_in_shift),
    .io_out_activate(PE_Array_14_24_io_out_activate),
    .io_out_weight(PE_Array_14_24_io_out_weight),
    .io_out_psum(PE_Array_14_24_io_out_psum)
  );
  basic_PE PE_Array_14_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_25_clock),
    .reset(PE_Array_14_25_reset),
    .io_in_activate(PE_Array_14_25_io_in_activate),
    .io_in_weight(PE_Array_14_25_io_in_weight),
    .io_in_psum(PE_Array_14_25_io_in_psum),
    .io_in_flow(PE_Array_14_25_io_in_flow),
    .io_in_shift(PE_Array_14_25_io_in_shift),
    .io_out_activate(PE_Array_14_25_io_out_activate),
    .io_out_weight(PE_Array_14_25_io_out_weight),
    .io_out_psum(PE_Array_14_25_io_out_psum)
  );
  basic_PE PE_Array_14_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_26_clock),
    .reset(PE_Array_14_26_reset),
    .io_in_activate(PE_Array_14_26_io_in_activate),
    .io_in_weight(PE_Array_14_26_io_in_weight),
    .io_in_psum(PE_Array_14_26_io_in_psum),
    .io_in_flow(PE_Array_14_26_io_in_flow),
    .io_in_shift(PE_Array_14_26_io_in_shift),
    .io_out_activate(PE_Array_14_26_io_out_activate),
    .io_out_weight(PE_Array_14_26_io_out_weight),
    .io_out_psum(PE_Array_14_26_io_out_psum)
  );
  basic_PE PE_Array_14_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_27_clock),
    .reset(PE_Array_14_27_reset),
    .io_in_activate(PE_Array_14_27_io_in_activate),
    .io_in_weight(PE_Array_14_27_io_in_weight),
    .io_in_psum(PE_Array_14_27_io_in_psum),
    .io_in_flow(PE_Array_14_27_io_in_flow),
    .io_in_shift(PE_Array_14_27_io_in_shift),
    .io_out_activate(PE_Array_14_27_io_out_activate),
    .io_out_weight(PE_Array_14_27_io_out_weight),
    .io_out_psum(PE_Array_14_27_io_out_psum)
  );
  basic_PE PE_Array_14_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_28_clock),
    .reset(PE_Array_14_28_reset),
    .io_in_activate(PE_Array_14_28_io_in_activate),
    .io_in_weight(PE_Array_14_28_io_in_weight),
    .io_in_psum(PE_Array_14_28_io_in_psum),
    .io_in_flow(PE_Array_14_28_io_in_flow),
    .io_in_shift(PE_Array_14_28_io_in_shift),
    .io_out_activate(PE_Array_14_28_io_out_activate),
    .io_out_weight(PE_Array_14_28_io_out_weight),
    .io_out_psum(PE_Array_14_28_io_out_psum)
  );
  basic_PE PE_Array_14_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_29_clock),
    .reset(PE_Array_14_29_reset),
    .io_in_activate(PE_Array_14_29_io_in_activate),
    .io_in_weight(PE_Array_14_29_io_in_weight),
    .io_in_psum(PE_Array_14_29_io_in_psum),
    .io_in_flow(PE_Array_14_29_io_in_flow),
    .io_in_shift(PE_Array_14_29_io_in_shift),
    .io_out_activate(PE_Array_14_29_io_out_activate),
    .io_out_weight(PE_Array_14_29_io_out_weight),
    .io_out_psum(PE_Array_14_29_io_out_psum)
  );
  basic_PE PE_Array_14_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_30_clock),
    .reset(PE_Array_14_30_reset),
    .io_in_activate(PE_Array_14_30_io_in_activate),
    .io_in_weight(PE_Array_14_30_io_in_weight),
    .io_in_psum(PE_Array_14_30_io_in_psum),
    .io_in_flow(PE_Array_14_30_io_in_flow),
    .io_in_shift(PE_Array_14_30_io_in_shift),
    .io_out_activate(PE_Array_14_30_io_out_activate),
    .io_out_weight(PE_Array_14_30_io_out_weight),
    .io_out_psum(PE_Array_14_30_io_out_psum)
  );
  basic_PE PE_Array_14_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_14_31_clock),
    .reset(PE_Array_14_31_reset),
    .io_in_activate(PE_Array_14_31_io_in_activate),
    .io_in_weight(PE_Array_14_31_io_in_weight),
    .io_in_psum(PE_Array_14_31_io_in_psum),
    .io_in_flow(PE_Array_14_31_io_in_flow),
    .io_in_shift(PE_Array_14_31_io_in_shift),
    .io_out_activate(PE_Array_14_31_io_out_activate),
    .io_out_weight(PE_Array_14_31_io_out_weight),
    .io_out_psum(PE_Array_14_31_io_out_psum)
  );
  basic_PE PE_Array_15_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_0_clock),
    .reset(PE_Array_15_0_reset),
    .io_in_activate(PE_Array_15_0_io_in_activate),
    .io_in_weight(PE_Array_15_0_io_in_weight),
    .io_in_psum(PE_Array_15_0_io_in_psum),
    .io_in_flow(PE_Array_15_0_io_in_flow),
    .io_in_shift(PE_Array_15_0_io_in_shift),
    .io_out_activate(PE_Array_15_0_io_out_activate),
    .io_out_weight(PE_Array_15_0_io_out_weight),
    .io_out_psum(PE_Array_15_0_io_out_psum)
  );
  basic_PE PE_Array_15_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_1_clock),
    .reset(PE_Array_15_1_reset),
    .io_in_activate(PE_Array_15_1_io_in_activate),
    .io_in_weight(PE_Array_15_1_io_in_weight),
    .io_in_psum(PE_Array_15_1_io_in_psum),
    .io_in_flow(PE_Array_15_1_io_in_flow),
    .io_in_shift(PE_Array_15_1_io_in_shift),
    .io_out_activate(PE_Array_15_1_io_out_activate),
    .io_out_weight(PE_Array_15_1_io_out_weight),
    .io_out_psum(PE_Array_15_1_io_out_psum)
  );
  basic_PE PE_Array_15_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_2_clock),
    .reset(PE_Array_15_2_reset),
    .io_in_activate(PE_Array_15_2_io_in_activate),
    .io_in_weight(PE_Array_15_2_io_in_weight),
    .io_in_psum(PE_Array_15_2_io_in_psum),
    .io_in_flow(PE_Array_15_2_io_in_flow),
    .io_in_shift(PE_Array_15_2_io_in_shift),
    .io_out_activate(PE_Array_15_2_io_out_activate),
    .io_out_weight(PE_Array_15_2_io_out_weight),
    .io_out_psum(PE_Array_15_2_io_out_psum)
  );
  basic_PE PE_Array_15_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_3_clock),
    .reset(PE_Array_15_3_reset),
    .io_in_activate(PE_Array_15_3_io_in_activate),
    .io_in_weight(PE_Array_15_3_io_in_weight),
    .io_in_psum(PE_Array_15_3_io_in_psum),
    .io_in_flow(PE_Array_15_3_io_in_flow),
    .io_in_shift(PE_Array_15_3_io_in_shift),
    .io_out_activate(PE_Array_15_3_io_out_activate),
    .io_out_weight(PE_Array_15_3_io_out_weight),
    .io_out_psum(PE_Array_15_3_io_out_psum)
  );
  basic_PE PE_Array_15_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_4_clock),
    .reset(PE_Array_15_4_reset),
    .io_in_activate(PE_Array_15_4_io_in_activate),
    .io_in_weight(PE_Array_15_4_io_in_weight),
    .io_in_psum(PE_Array_15_4_io_in_psum),
    .io_in_flow(PE_Array_15_4_io_in_flow),
    .io_in_shift(PE_Array_15_4_io_in_shift),
    .io_out_activate(PE_Array_15_4_io_out_activate),
    .io_out_weight(PE_Array_15_4_io_out_weight),
    .io_out_psum(PE_Array_15_4_io_out_psum)
  );
  basic_PE PE_Array_15_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_5_clock),
    .reset(PE_Array_15_5_reset),
    .io_in_activate(PE_Array_15_5_io_in_activate),
    .io_in_weight(PE_Array_15_5_io_in_weight),
    .io_in_psum(PE_Array_15_5_io_in_psum),
    .io_in_flow(PE_Array_15_5_io_in_flow),
    .io_in_shift(PE_Array_15_5_io_in_shift),
    .io_out_activate(PE_Array_15_5_io_out_activate),
    .io_out_weight(PE_Array_15_5_io_out_weight),
    .io_out_psum(PE_Array_15_5_io_out_psum)
  );
  basic_PE PE_Array_15_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_6_clock),
    .reset(PE_Array_15_6_reset),
    .io_in_activate(PE_Array_15_6_io_in_activate),
    .io_in_weight(PE_Array_15_6_io_in_weight),
    .io_in_psum(PE_Array_15_6_io_in_psum),
    .io_in_flow(PE_Array_15_6_io_in_flow),
    .io_in_shift(PE_Array_15_6_io_in_shift),
    .io_out_activate(PE_Array_15_6_io_out_activate),
    .io_out_weight(PE_Array_15_6_io_out_weight),
    .io_out_psum(PE_Array_15_6_io_out_psum)
  );
  basic_PE PE_Array_15_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_7_clock),
    .reset(PE_Array_15_7_reset),
    .io_in_activate(PE_Array_15_7_io_in_activate),
    .io_in_weight(PE_Array_15_7_io_in_weight),
    .io_in_psum(PE_Array_15_7_io_in_psum),
    .io_in_flow(PE_Array_15_7_io_in_flow),
    .io_in_shift(PE_Array_15_7_io_in_shift),
    .io_out_activate(PE_Array_15_7_io_out_activate),
    .io_out_weight(PE_Array_15_7_io_out_weight),
    .io_out_psum(PE_Array_15_7_io_out_psum)
  );
  basic_PE PE_Array_15_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_8_clock),
    .reset(PE_Array_15_8_reset),
    .io_in_activate(PE_Array_15_8_io_in_activate),
    .io_in_weight(PE_Array_15_8_io_in_weight),
    .io_in_psum(PE_Array_15_8_io_in_psum),
    .io_in_flow(PE_Array_15_8_io_in_flow),
    .io_in_shift(PE_Array_15_8_io_in_shift),
    .io_out_activate(PE_Array_15_8_io_out_activate),
    .io_out_weight(PE_Array_15_8_io_out_weight),
    .io_out_psum(PE_Array_15_8_io_out_psum)
  );
  basic_PE PE_Array_15_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_9_clock),
    .reset(PE_Array_15_9_reset),
    .io_in_activate(PE_Array_15_9_io_in_activate),
    .io_in_weight(PE_Array_15_9_io_in_weight),
    .io_in_psum(PE_Array_15_9_io_in_psum),
    .io_in_flow(PE_Array_15_9_io_in_flow),
    .io_in_shift(PE_Array_15_9_io_in_shift),
    .io_out_activate(PE_Array_15_9_io_out_activate),
    .io_out_weight(PE_Array_15_9_io_out_weight),
    .io_out_psum(PE_Array_15_9_io_out_psum)
  );
  basic_PE PE_Array_15_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_10_clock),
    .reset(PE_Array_15_10_reset),
    .io_in_activate(PE_Array_15_10_io_in_activate),
    .io_in_weight(PE_Array_15_10_io_in_weight),
    .io_in_psum(PE_Array_15_10_io_in_psum),
    .io_in_flow(PE_Array_15_10_io_in_flow),
    .io_in_shift(PE_Array_15_10_io_in_shift),
    .io_out_activate(PE_Array_15_10_io_out_activate),
    .io_out_weight(PE_Array_15_10_io_out_weight),
    .io_out_psum(PE_Array_15_10_io_out_psum)
  );
  basic_PE PE_Array_15_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_11_clock),
    .reset(PE_Array_15_11_reset),
    .io_in_activate(PE_Array_15_11_io_in_activate),
    .io_in_weight(PE_Array_15_11_io_in_weight),
    .io_in_psum(PE_Array_15_11_io_in_psum),
    .io_in_flow(PE_Array_15_11_io_in_flow),
    .io_in_shift(PE_Array_15_11_io_in_shift),
    .io_out_activate(PE_Array_15_11_io_out_activate),
    .io_out_weight(PE_Array_15_11_io_out_weight),
    .io_out_psum(PE_Array_15_11_io_out_psum)
  );
  basic_PE PE_Array_15_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_12_clock),
    .reset(PE_Array_15_12_reset),
    .io_in_activate(PE_Array_15_12_io_in_activate),
    .io_in_weight(PE_Array_15_12_io_in_weight),
    .io_in_psum(PE_Array_15_12_io_in_psum),
    .io_in_flow(PE_Array_15_12_io_in_flow),
    .io_in_shift(PE_Array_15_12_io_in_shift),
    .io_out_activate(PE_Array_15_12_io_out_activate),
    .io_out_weight(PE_Array_15_12_io_out_weight),
    .io_out_psum(PE_Array_15_12_io_out_psum)
  );
  basic_PE PE_Array_15_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_13_clock),
    .reset(PE_Array_15_13_reset),
    .io_in_activate(PE_Array_15_13_io_in_activate),
    .io_in_weight(PE_Array_15_13_io_in_weight),
    .io_in_psum(PE_Array_15_13_io_in_psum),
    .io_in_flow(PE_Array_15_13_io_in_flow),
    .io_in_shift(PE_Array_15_13_io_in_shift),
    .io_out_activate(PE_Array_15_13_io_out_activate),
    .io_out_weight(PE_Array_15_13_io_out_weight),
    .io_out_psum(PE_Array_15_13_io_out_psum)
  );
  basic_PE PE_Array_15_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_14_clock),
    .reset(PE_Array_15_14_reset),
    .io_in_activate(PE_Array_15_14_io_in_activate),
    .io_in_weight(PE_Array_15_14_io_in_weight),
    .io_in_psum(PE_Array_15_14_io_in_psum),
    .io_in_flow(PE_Array_15_14_io_in_flow),
    .io_in_shift(PE_Array_15_14_io_in_shift),
    .io_out_activate(PE_Array_15_14_io_out_activate),
    .io_out_weight(PE_Array_15_14_io_out_weight),
    .io_out_psum(PE_Array_15_14_io_out_psum)
  );
  basic_PE PE_Array_15_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_15_clock),
    .reset(PE_Array_15_15_reset),
    .io_in_activate(PE_Array_15_15_io_in_activate),
    .io_in_weight(PE_Array_15_15_io_in_weight),
    .io_in_psum(PE_Array_15_15_io_in_psum),
    .io_in_flow(PE_Array_15_15_io_in_flow),
    .io_in_shift(PE_Array_15_15_io_in_shift),
    .io_out_activate(PE_Array_15_15_io_out_activate),
    .io_out_weight(PE_Array_15_15_io_out_weight),
    .io_out_psum(PE_Array_15_15_io_out_psum)
  );
  basic_PE PE_Array_15_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_16_clock),
    .reset(PE_Array_15_16_reset),
    .io_in_activate(PE_Array_15_16_io_in_activate),
    .io_in_weight(PE_Array_15_16_io_in_weight),
    .io_in_psum(PE_Array_15_16_io_in_psum),
    .io_in_flow(PE_Array_15_16_io_in_flow),
    .io_in_shift(PE_Array_15_16_io_in_shift),
    .io_out_activate(PE_Array_15_16_io_out_activate),
    .io_out_weight(PE_Array_15_16_io_out_weight),
    .io_out_psum(PE_Array_15_16_io_out_psum)
  );
  basic_PE PE_Array_15_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_17_clock),
    .reset(PE_Array_15_17_reset),
    .io_in_activate(PE_Array_15_17_io_in_activate),
    .io_in_weight(PE_Array_15_17_io_in_weight),
    .io_in_psum(PE_Array_15_17_io_in_psum),
    .io_in_flow(PE_Array_15_17_io_in_flow),
    .io_in_shift(PE_Array_15_17_io_in_shift),
    .io_out_activate(PE_Array_15_17_io_out_activate),
    .io_out_weight(PE_Array_15_17_io_out_weight),
    .io_out_psum(PE_Array_15_17_io_out_psum)
  );
  basic_PE PE_Array_15_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_18_clock),
    .reset(PE_Array_15_18_reset),
    .io_in_activate(PE_Array_15_18_io_in_activate),
    .io_in_weight(PE_Array_15_18_io_in_weight),
    .io_in_psum(PE_Array_15_18_io_in_psum),
    .io_in_flow(PE_Array_15_18_io_in_flow),
    .io_in_shift(PE_Array_15_18_io_in_shift),
    .io_out_activate(PE_Array_15_18_io_out_activate),
    .io_out_weight(PE_Array_15_18_io_out_weight),
    .io_out_psum(PE_Array_15_18_io_out_psum)
  );
  basic_PE PE_Array_15_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_19_clock),
    .reset(PE_Array_15_19_reset),
    .io_in_activate(PE_Array_15_19_io_in_activate),
    .io_in_weight(PE_Array_15_19_io_in_weight),
    .io_in_psum(PE_Array_15_19_io_in_psum),
    .io_in_flow(PE_Array_15_19_io_in_flow),
    .io_in_shift(PE_Array_15_19_io_in_shift),
    .io_out_activate(PE_Array_15_19_io_out_activate),
    .io_out_weight(PE_Array_15_19_io_out_weight),
    .io_out_psum(PE_Array_15_19_io_out_psum)
  );
  basic_PE PE_Array_15_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_20_clock),
    .reset(PE_Array_15_20_reset),
    .io_in_activate(PE_Array_15_20_io_in_activate),
    .io_in_weight(PE_Array_15_20_io_in_weight),
    .io_in_psum(PE_Array_15_20_io_in_psum),
    .io_in_flow(PE_Array_15_20_io_in_flow),
    .io_in_shift(PE_Array_15_20_io_in_shift),
    .io_out_activate(PE_Array_15_20_io_out_activate),
    .io_out_weight(PE_Array_15_20_io_out_weight),
    .io_out_psum(PE_Array_15_20_io_out_psum)
  );
  basic_PE PE_Array_15_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_21_clock),
    .reset(PE_Array_15_21_reset),
    .io_in_activate(PE_Array_15_21_io_in_activate),
    .io_in_weight(PE_Array_15_21_io_in_weight),
    .io_in_psum(PE_Array_15_21_io_in_psum),
    .io_in_flow(PE_Array_15_21_io_in_flow),
    .io_in_shift(PE_Array_15_21_io_in_shift),
    .io_out_activate(PE_Array_15_21_io_out_activate),
    .io_out_weight(PE_Array_15_21_io_out_weight),
    .io_out_psum(PE_Array_15_21_io_out_psum)
  );
  basic_PE PE_Array_15_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_22_clock),
    .reset(PE_Array_15_22_reset),
    .io_in_activate(PE_Array_15_22_io_in_activate),
    .io_in_weight(PE_Array_15_22_io_in_weight),
    .io_in_psum(PE_Array_15_22_io_in_psum),
    .io_in_flow(PE_Array_15_22_io_in_flow),
    .io_in_shift(PE_Array_15_22_io_in_shift),
    .io_out_activate(PE_Array_15_22_io_out_activate),
    .io_out_weight(PE_Array_15_22_io_out_weight),
    .io_out_psum(PE_Array_15_22_io_out_psum)
  );
  basic_PE PE_Array_15_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_23_clock),
    .reset(PE_Array_15_23_reset),
    .io_in_activate(PE_Array_15_23_io_in_activate),
    .io_in_weight(PE_Array_15_23_io_in_weight),
    .io_in_psum(PE_Array_15_23_io_in_psum),
    .io_in_flow(PE_Array_15_23_io_in_flow),
    .io_in_shift(PE_Array_15_23_io_in_shift),
    .io_out_activate(PE_Array_15_23_io_out_activate),
    .io_out_weight(PE_Array_15_23_io_out_weight),
    .io_out_psum(PE_Array_15_23_io_out_psum)
  );
  basic_PE PE_Array_15_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_24_clock),
    .reset(PE_Array_15_24_reset),
    .io_in_activate(PE_Array_15_24_io_in_activate),
    .io_in_weight(PE_Array_15_24_io_in_weight),
    .io_in_psum(PE_Array_15_24_io_in_psum),
    .io_in_flow(PE_Array_15_24_io_in_flow),
    .io_in_shift(PE_Array_15_24_io_in_shift),
    .io_out_activate(PE_Array_15_24_io_out_activate),
    .io_out_weight(PE_Array_15_24_io_out_weight),
    .io_out_psum(PE_Array_15_24_io_out_psum)
  );
  basic_PE PE_Array_15_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_25_clock),
    .reset(PE_Array_15_25_reset),
    .io_in_activate(PE_Array_15_25_io_in_activate),
    .io_in_weight(PE_Array_15_25_io_in_weight),
    .io_in_psum(PE_Array_15_25_io_in_psum),
    .io_in_flow(PE_Array_15_25_io_in_flow),
    .io_in_shift(PE_Array_15_25_io_in_shift),
    .io_out_activate(PE_Array_15_25_io_out_activate),
    .io_out_weight(PE_Array_15_25_io_out_weight),
    .io_out_psum(PE_Array_15_25_io_out_psum)
  );
  basic_PE PE_Array_15_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_26_clock),
    .reset(PE_Array_15_26_reset),
    .io_in_activate(PE_Array_15_26_io_in_activate),
    .io_in_weight(PE_Array_15_26_io_in_weight),
    .io_in_psum(PE_Array_15_26_io_in_psum),
    .io_in_flow(PE_Array_15_26_io_in_flow),
    .io_in_shift(PE_Array_15_26_io_in_shift),
    .io_out_activate(PE_Array_15_26_io_out_activate),
    .io_out_weight(PE_Array_15_26_io_out_weight),
    .io_out_psum(PE_Array_15_26_io_out_psum)
  );
  basic_PE PE_Array_15_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_27_clock),
    .reset(PE_Array_15_27_reset),
    .io_in_activate(PE_Array_15_27_io_in_activate),
    .io_in_weight(PE_Array_15_27_io_in_weight),
    .io_in_psum(PE_Array_15_27_io_in_psum),
    .io_in_flow(PE_Array_15_27_io_in_flow),
    .io_in_shift(PE_Array_15_27_io_in_shift),
    .io_out_activate(PE_Array_15_27_io_out_activate),
    .io_out_weight(PE_Array_15_27_io_out_weight),
    .io_out_psum(PE_Array_15_27_io_out_psum)
  );
  basic_PE PE_Array_15_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_28_clock),
    .reset(PE_Array_15_28_reset),
    .io_in_activate(PE_Array_15_28_io_in_activate),
    .io_in_weight(PE_Array_15_28_io_in_weight),
    .io_in_psum(PE_Array_15_28_io_in_psum),
    .io_in_flow(PE_Array_15_28_io_in_flow),
    .io_in_shift(PE_Array_15_28_io_in_shift),
    .io_out_activate(PE_Array_15_28_io_out_activate),
    .io_out_weight(PE_Array_15_28_io_out_weight),
    .io_out_psum(PE_Array_15_28_io_out_psum)
  );
  basic_PE PE_Array_15_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_29_clock),
    .reset(PE_Array_15_29_reset),
    .io_in_activate(PE_Array_15_29_io_in_activate),
    .io_in_weight(PE_Array_15_29_io_in_weight),
    .io_in_psum(PE_Array_15_29_io_in_psum),
    .io_in_flow(PE_Array_15_29_io_in_flow),
    .io_in_shift(PE_Array_15_29_io_in_shift),
    .io_out_activate(PE_Array_15_29_io_out_activate),
    .io_out_weight(PE_Array_15_29_io_out_weight),
    .io_out_psum(PE_Array_15_29_io_out_psum)
  );
  basic_PE PE_Array_15_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_30_clock),
    .reset(PE_Array_15_30_reset),
    .io_in_activate(PE_Array_15_30_io_in_activate),
    .io_in_weight(PE_Array_15_30_io_in_weight),
    .io_in_psum(PE_Array_15_30_io_in_psum),
    .io_in_flow(PE_Array_15_30_io_in_flow),
    .io_in_shift(PE_Array_15_30_io_in_shift),
    .io_out_activate(PE_Array_15_30_io_out_activate),
    .io_out_weight(PE_Array_15_30_io_out_weight),
    .io_out_psum(PE_Array_15_30_io_out_psum)
  );
  basic_PE PE_Array_15_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_15_31_clock),
    .reset(PE_Array_15_31_reset),
    .io_in_activate(PE_Array_15_31_io_in_activate),
    .io_in_weight(PE_Array_15_31_io_in_weight),
    .io_in_psum(PE_Array_15_31_io_in_psum),
    .io_in_flow(PE_Array_15_31_io_in_flow),
    .io_in_shift(PE_Array_15_31_io_in_shift),
    .io_out_activate(PE_Array_15_31_io_out_activate),
    .io_out_weight(PE_Array_15_31_io_out_weight),
    .io_out_psum(PE_Array_15_31_io_out_psum)
  );
  basic_PE PE_Array_16_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_0_clock),
    .reset(PE_Array_16_0_reset),
    .io_in_activate(PE_Array_16_0_io_in_activate),
    .io_in_weight(PE_Array_16_0_io_in_weight),
    .io_in_psum(PE_Array_16_0_io_in_psum),
    .io_in_flow(PE_Array_16_0_io_in_flow),
    .io_in_shift(PE_Array_16_0_io_in_shift),
    .io_out_activate(PE_Array_16_0_io_out_activate),
    .io_out_weight(PE_Array_16_0_io_out_weight),
    .io_out_psum(PE_Array_16_0_io_out_psum)
  );
  basic_PE PE_Array_16_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_1_clock),
    .reset(PE_Array_16_1_reset),
    .io_in_activate(PE_Array_16_1_io_in_activate),
    .io_in_weight(PE_Array_16_1_io_in_weight),
    .io_in_psum(PE_Array_16_1_io_in_psum),
    .io_in_flow(PE_Array_16_1_io_in_flow),
    .io_in_shift(PE_Array_16_1_io_in_shift),
    .io_out_activate(PE_Array_16_1_io_out_activate),
    .io_out_weight(PE_Array_16_1_io_out_weight),
    .io_out_psum(PE_Array_16_1_io_out_psum)
  );
  basic_PE PE_Array_16_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_2_clock),
    .reset(PE_Array_16_2_reset),
    .io_in_activate(PE_Array_16_2_io_in_activate),
    .io_in_weight(PE_Array_16_2_io_in_weight),
    .io_in_psum(PE_Array_16_2_io_in_psum),
    .io_in_flow(PE_Array_16_2_io_in_flow),
    .io_in_shift(PE_Array_16_2_io_in_shift),
    .io_out_activate(PE_Array_16_2_io_out_activate),
    .io_out_weight(PE_Array_16_2_io_out_weight),
    .io_out_psum(PE_Array_16_2_io_out_psum)
  );
  basic_PE PE_Array_16_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_3_clock),
    .reset(PE_Array_16_3_reset),
    .io_in_activate(PE_Array_16_3_io_in_activate),
    .io_in_weight(PE_Array_16_3_io_in_weight),
    .io_in_psum(PE_Array_16_3_io_in_psum),
    .io_in_flow(PE_Array_16_3_io_in_flow),
    .io_in_shift(PE_Array_16_3_io_in_shift),
    .io_out_activate(PE_Array_16_3_io_out_activate),
    .io_out_weight(PE_Array_16_3_io_out_weight),
    .io_out_psum(PE_Array_16_3_io_out_psum)
  );
  basic_PE PE_Array_16_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_4_clock),
    .reset(PE_Array_16_4_reset),
    .io_in_activate(PE_Array_16_4_io_in_activate),
    .io_in_weight(PE_Array_16_4_io_in_weight),
    .io_in_psum(PE_Array_16_4_io_in_psum),
    .io_in_flow(PE_Array_16_4_io_in_flow),
    .io_in_shift(PE_Array_16_4_io_in_shift),
    .io_out_activate(PE_Array_16_4_io_out_activate),
    .io_out_weight(PE_Array_16_4_io_out_weight),
    .io_out_psum(PE_Array_16_4_io_out_psum)
  );
  basic_PE PE_Array_16_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_5_clock),
    .reset(PE_Array_16_5_reset),
    .io_in_activate(PE_Array_16_5_io_in_activate),
    .io_in_weight(PE_Array_16_5_io_in_weight),
    .io_in_psum(PE_Array_16_5_io_in_psum),
    .io_in_flow(PE_Array_16_5_io_in_flow),
    .io_in_shift(PE_Array_16_5_io_in_shift),
    .io_out_activate(PE_Array_16_5_io_out_activate),
    .io_out_weight(PE_Array_16_5_io_out_weight),
    .io_out_psum(PE_Array_16_5_io_out_psum)
  );
  basic_PE PE_Array_16_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_6_clock),
    .reset(PE_Array_16_6_reset),
    .io_in_activate(PE_Array_16_6_io_in_activate),
    .io_in_weight(PE_Array_16_6_io_in_weight),
    .io_in_psum(PE_Array_16_6_io_in_psum),
    .io_in_flow(PE_Array_16_6_io_in_flow),
    .io_in_shift(PE_Array_16_6_io_in_shift),
    .io_out_activate(PE_Array_16_6_io_out_activate),
    .io_out_weight(PE_Array_16_6_io_out_weight),
    .io_out_psum(PE_Array_16_6_io_out_psum)
  );
  basic_PE PE_Array_16_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_7_clock),
    .reset(PE_Array_16_7_reset),
    .io_in_activate(PE_Array_16_7_io_in_activate),
    .io_in_weight(PE_Array_16_7_io_in_weight),
    .io_in_psum(PE_Array_16_7_io_in_psum),
    .io_in_flow(PE_Array_16_7_io_in_flow),
    .io_in_shift(PE_Array_16_7_io_in_shift),
    .io_out_activate(PE_Array_16_7_io_out_activate),
    .io_out_weight(PE_Array_16_7_io_out_weight),
    .io_out_psum(PE_Array_16_7_io_out_psum)
  );
  basic_PE PE_Array_16_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_8_clock),
    .reset(PE_Array_16_8_reset),
    .io_in_activate(PE_Array_16_8_io_in_activate),
    .io_in_weight(PE_Array_16_8_io_in_weight),
    .io_in_psum(PE_Array_16_8_io_in_psum),
    .io_in_flow(PE_Array_16_8_io_in_flow),
    .io_in_shift(PE_Array_16_8_io_in_shift),
    .io_out_activate(PE_Array_16_8_io_out_activate),
    .io_out_weight(PE_Array_16_8_io_out_weight),
    .io_out_psum(PE_Array_16_8_io_out_psum)
  );
  basic_PE PE_Array_16_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_9_clock),
    .reset(PE_Array_16_9_reset),
    .io_in_activate(PE_Array_16_9_io_in_activate),
    .io_in_weight(PE_Array_16_9_io_in_weight),
    .io_in_psum(PE_Array_16_9_io_in_psum),
    .io_in_flow(PE_Array_16_9_io_in_flow),
    .io_in_shift(PE_Array_16_9_io_in_shift),
    .io_out_activate(PE_Array_16_9_io_out_activate),
    .io_out_weight(PE_Array_16_9_io_out_weight),
    .io_out_psum(PE_Array_16_9_io_out_psum)
  );
  basic_PE PE_Array_16_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_10_clock),
    .reset(PE_Array_16_10_reset),
    .io_in_activate(PE_Array_16_10_io_in_activate),
    .io_in_weight(PE_Array_16_10_io_in_weight),
    .io_in_psum(PE_Array_16_10_io_in_psum),
    .io_in_flow(PE_Array_16_10_io_in_flow),
    .io_in_shift(PE_Array_16_10_io_in_shift),
    .io_out_activate(PE_Array_16_10_io_out_activate),
    .io_out_weight(PE_Array_16_10_io_out_weight),
    .io_out_psum(PE_Array_16_10_io_out_psum)
  );
  basic_PE PE_Array_16_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_11_clock),
    .reset(PE_Array_16_11_reset),
    .io_in_activate(PE_Array_16_11_io_in_activate),
    .io_in_weight(PE_Array_16_11_io_in_weight),
    .io_in_psum(PE_Array_16_11_io_in_psum),
    .io_in_flow(PE_Array_16_11_io_in_flow),
    .io_in_shift(PE_Array_16_11_io_in_shift),
    .io_out_activate(PE_Array_16_11_io_out_activate),
    .io_out_weight(PE_Array_16_11_io_out_weight),
    .io_out_psum(PE_Array_16_11_io_out_psum)
  );
  basic_PE PE_Array_16_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_12_clock),
    .reset(PE_Array_16_12_reset),
    .io_in_activate(PE_Array_16_12_io_in_activate),
    .io_in_weight(PE_Array_16_12_io_in_weight),
    .io_in_psum(PE_Array_16_12_io_in_psum),
    .io_in_flow(PE_Array_16_12_io_in_flow),
    .io_in_shift(PE_Array_16_12_io_in_shift),
    .io_out_activate(PE_Array_16_12_io_out_activate),
    .io_out_weight(PE_Array_16_12_io_out_weight),
    .io_out_psum(PE_Array_16_12_io_out_psum)
  );
  basic_PE PE_Array_16_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_13_clock),
    .reset(PE_Array_16_13_reset),
    .io_in_activate(PE_Array_16_13_io_in_activate),
    .io_in_weight(PE_Array_16_13_io_in_weight),
    .io_in_psum(PE_Array_16_13_io_in_psum),
    .io_in_flow(PE_Array_16_13_io_in_flow),
    .io_in_shift(PE_Array_16_13_io_in_shift),
    .io_out_activate(PE_Array_16_13_io_out_activate),
    .io_out_weight(PE_Array_16_13_io_out_weight),
    .io_out_psum(PE_Array_16_13_io_out_psum)
  );
  basic_PE PE_Array_16_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_14_clock),
    .reset(PE_Array_16_14_reset),
    .io_in_activate(PE_Array_16_14_io_in_activate),
    .io_in_weight(PE_Array_16_14_io_in_weight),
    .io_in_psum(PE_Array_16_14_io_in_psum),
    .io_in_flow(PE_Array_16_14_io_in_flow),
    .io_in_shift(PE_Array_16_14_io_in_shift),
    .io_out_activate(PE_Array_16_14_io_out_activate),
    .io_out_weight(PE_Array_16_14_io_out_weight),
    .io_out_psum(PE_Array_16_14_io_out_psum)
  );
  basic_PE PE_Array_16_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_15_clock),
    .reset(PE_Array_16_15_reset),
    .io_in_activate(PE_Array_16_15_io_in_activate),
    .io_in_weight(PE_Array_16_15_io_in_weight),
    .io_in_psum(PE_Array_16_15_io_in_psum),
    .io_in_flow(PE_Array_16_15_io_in_flow),
    .io_in_shift(PE_Array_16_15_io_in_shift),
    .io_out_activate(PE_Array_16_15_io_out_activate),
    .io_out_weight(PE_Array_16_15_io_out_weight),
    .io_out_psum(PE_Array_16_15_io_out_psum)
  );
  basic_PE PE_Array_16_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_16_clock),
    .reset(PE_Array_16_16_reset),
    .io_in_activate(PE_Array_16_16_io_in_activate),
    .io_in_weight(PE_Array_16_16_io_in_weight),
    .io_in_psum(PE_Array_16_16_io_in_psum),
    .io_in_flow(PE_Array_16_16_io_in_flow),
    .io_in_shift(PE_Array_16_16_io_in_shift),
    .io_out_activate(PE_Array_16_16_io_out_activate),
    .io_out_weight(PE_Array_16_16_io_out_weight),
    .io_out_psum(PE_Array_16_16_io_out_psum)
  );
  basic_PE PE_Array_16_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_17_clock),
    .reset(PE_Array_16_17_reset),
    .io_in_activate(PE_Array_16_17_io_in_activate),
    .io_in_weight(PE_Array_16_17_io_in_weight),
    .io_in_psum(PE_Array_16_17_io_in_psum),
    .io_in_flow(PE_Array_16_17_io_in_flow),
    .io_in_shift(PE_Array_16_17_io_in_shift),
    .io_out_activate(PE_Array_16_17_io_out_activate),
    .io_out_weight(PE_Array_16_17_io_out_weight),
    .io_out_psum(PE_Array_16_17_io_out_psum)
  );
  basic_PE PE_Array_16_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_18_clock),
    .reset(PE_Array_16_18_reset),
    .io_in_activate(PE_Array_16_18_io_in_activate),
    .io_in_weight(PE_Array_16_18_io_in_weight),
    .io_in_psum(PE_Array_16_18_io_in_psum),
    .io_in_flow(PE_Array_16_18_io_in_flow),
    .io_in_shift(PE_Array_16_18_io_in_shift),
    .io_out_activate(PE_Array_16_18_io_out_activate),
    .io_out_weight(PE_Array_16_18_io_out_weight),
    .io_out_psum(PE_Array_16_18_io_out_psum)
  );
  basic_PE PE_Array_16_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_19_clock),
    .reset(PE_Array_16_19_reset),
    .io_in_activate(PE_Array_16_19_io_in_activate),
    .io_in_weight(PE_Array_16_19_io_in_weight),
    .io_in_psum(PE_Array_16_19_io_in_psum),
    .io_in_flow(PE_Array_16_19_io_in_flow),
    .io_in_shift(PE_Array_16_19_io_in_shift),
    .io_out_activate(PE_Array_16_19_io_out_activate),
    .io_out_weight(PE_Array_16_19_io_out_weight),
    .io_out_psum(PE_Array_16_19_io_out_psum)
  );
  basic_PE PE_Array_16_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_20_clock),
    .reset(PE_Array_16_20_reset),
    .io_in_activate(PE_Array_16_20_io_in_activate),
    .io_in_weight(PE_Array_16_20_io_in_weight),
    .io_in_psum(PE_Array_16_20_io_in_psum),
    .io_in_flow(PE_Array_16_20_io_in_flow),
    .io_in_shift(PE_Array_16_20_io_in_shift),
    .io_out_activate(PE_Array_16_20_io_out_activate),
    .io_out_weight(PE_Array_16_20_io_out_weight),
    .io_out_psum(PE_Array_16_20_io_out_psum)
  );
  basic_PE PE_Array_16_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_21_clock),
    .reset(PE_Array_16_21_reset),
    .io_in_activate(PE_Array_16_21_io_in_activate),
    .io_in_weight(PE_Array_16_21_io_in_weight),
    .io_in_psum(PE_Array_16_21_io_in_psum),
    .io_in_flow(PE_Array_16_21_io_in_flow),
    .io_in_shift(PE_Array_16_21_io_in_shift),
    .io_out_activate(PE_Array_16_21_io_out_activate),
    .io_out_weight(PE_Array_16_21_io_out_weight),
    .io_out_psum(PE_Array_16_21_io_out_psum)
  );
  basic_PE PE_Array_16_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_22_clock),
    .reset(PE_Array_16_22_reset),
    .io_in_activate(PE_Array_16_22_io_in_activate),
    .io_in_weight(PE_Array_16_22_io_in_weight),
    .io_in_psum(PE_Array_16_22_io_in_psum),
    .io_in_flow(PE_Array_16_22_io_in_flow),
    .io_in_shift(PE_Array_16_22_io_in_shift),
    .io_out_activate(PE_Array_16_22_io_out_activate),
    .io_out_weight(PE_Array_16_22_io_out_weight),
    .io_out_psum(PE_Array_16_22_io_out_psum)
  );
  basic_PE PE_Array_16_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_23_clock),
    .reset(PE_Array_16_23_reset),
    .io_in_activate(PE_Array_16_23_io_in_activate),
    .io_in_weight(PE_Array_16_23_io_in_weight),
    .io_in_psum(PE_Array_16_23_io_in_psum),
    .io_in_flow(PE_Array_16_23_io_in_flow),
    .io_in_shift(PE_Array_16_23_io_in_shift),
    .io_out_activate(PE_Array_16_23_io_out_activate),
    .io_out_weight(PE_Array_16_23_io_out_weight),
    .io_out_psum(PE_Array_16_23_io_out_psum)
  );
  basic_PE PE_Array_16_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_24_clock),
    .reset(PE_Array_16_24_reset),
    .io_in_activate(PE_Array_16_24_io_in_activate),
    .io_in_weight(PE_Array_16_24_io_in_weight),
    .io_in_psum(PE_Array_16_24_io_in_psum),
    .io_in_flow(PE_Array_16_24_io_in_flow),
    .io_in_shift(PE_Array_16_24_io_in_shift),
    .io_out_activate(PE_Array_16_24_io_out_activate),
    .io_out_weight(PE_Array_16_24_io_out_weight),
    .io_out_psum(PE_Array_16_24_io_out_psum)
  );
  basic_PE PE_Array_16_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_25_clock),
    .reset(PE_Array_16_25_reset),
    .io_in_activate(PE_Array_16_25_io_in_activate),
    .io_in_weight(PE_Array_16_25_io_in_weight),
    .io_in_psum(PE_Array_16_25_io_in_psum),
    .io_in_flow(PE_Array_16_25_io_in_flow),
    .io_in_shift(PE_Array_16_25_io_in_shift),
    .io_out_activate(PE_Array_16_25_io_out_activate),
    .io_out_weight(PE_Array_16_25_io_out_weight),
    .io_out_psum(PE_Array_16_25_io_out_psum)
  );
  basic_PE PE_Array_16_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_26_clock),
    .reset(PE_Array_16_26_reset),
    .io_in_activate(PE_Array_16_26_io_in_activate),
    .io_in_weight(PE_Array_16_26_io_in_weight),
    .io_in_psum(PE_Array_16_26_io_in_psum),
    .io_in_flow(PE_Array_16_26_io_in_flow),
    .io_in_shift(PE_Array_16_26_io_in_shift),
    .io_out_activate(PE_Array_16_26_io_out_activate),
    .io_out_weight(PE_Array_16_26_io_out_weight),
    .io_out_psum(PE_Array_16_26_io_out_psum)
  );
  basic_PE PE_Array_16_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_27_clock),
    .reset(PE_Array_16_27_reset),
    .io_in_activate(PE_Array_16_27_io_in_activate),
    .io_in_weight(PE_Array_16_27_io_in_weight),
    .io_in_psum(PE_Array_16_27_io_in_psum),
    .io_in_flow(PE_Array_16_27_io_in_flow),
    .io_in_shift(PE_Array_16_27_io_in_shift),
    .io_out_activate(PE_Array_16_27_io_out_activate),
    .io_out_weight(PE_Array_16_27_io_out_weight),
    .io_out_psum(PE_Array_16_27_io_out_psum)
  );
  basic_PE PE_Array_16_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_28_clock),
    .reset(PE_Array_16_28_reset),
    .io_in_activate(PE_Array_16_28_io_in_activate),
    .io_in_weight(PE_Array_16_28_io_in_weight),
    .io_in_psum(PE_Array_16_28_io_in_psum),
    .io_in_flow(PE_Array_16_28_io_in_flow),
    .io_in_shift(PE_Array_16_28_io_in_shift),
    .io_out_activate(PE_Array_16_28_io_out_activate),
    .io_out_weight(PE_Array_16_28_io_out_weight),
    .io_out_psum(PE_Array_16_28_io_out_psum)
  );
  basic_PE PE_Array_16_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_29_clock),
    .reset(PE_Array_16_29_reset),
    .io_in_activate(PE_Array_16_29_io_in_activate),
    .io_in_weight(PE_Array_16_29_io_in_weight),
    .io_in_psum(PE_Array_16_29_io_in_psum),
    .io_in_flow(PE_Array_16_29_io_in_flow),
    .io_in_shift(PE_Array_16_29_io_in_shift),
    .io_out_activate(PE_Array_16_29_io_out_activate),
    .io_out_weight(PE_Array_16_29_io_out_weight),
    .io_out_psum(PE_Array_16_29_io_out_psum)
  );
  basic_PE PE_Array_16_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_30_clock),
    .reset(PE_Array_16_30_reset),
    .io_in_activate(PE_Array_16_30_io_in_activate),
    .io_in_weight(PE_Array_16_30_io_in_weight),
    .io_in_psum(PE_Array_16_30_io_in_psum),
    .io_in_flow(PE_Array_16_30_io_in_flow),
    .io_in_shift(PE_Array_16_30_io_in_shift),
    .io_out_activate(PE_Array_16_30_io_out_activate),
    .io_out_weight(PE_Array_16_30_io_out_weight),
    .io_out_psum(PE_Array_16_30_io_out_psum)
  );
  basic_PE PE_Array_16_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_16_31_clock),
    .reset(PE_Array_16_31_reset),
    .io_in_activate(PE_Array_16_31_io_in_activate),
    .io_in_weight(PE_Array_16_31_io_in_weight),
    .io_in_psum(PE_Array_16_31_io_in_psum),
    .io_in_flow(PE_Array_16_31_io_in_flow),
    .io_in_shift(PE_Array_16_31_io_in_shift),
    .io_out_activate(PE_Array_16_31_io_out_activate),
    .io_out_weight(PE_Array_16_31_io_out_weight),
    .io_out_psum(PE_Array_16_31_io_out_psum)
  );
  basic_PE PE_Array_17_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_0_clock),
    .reset(PE_Array_17_0_reset),
    .io_in_activate(PE_Array_17_0_io_in_activate),
    .io_in_weight(PE_Array_17_0_io_in_weight),
    .io_in_psum(PE_Array_17_0_io_in_psum),
    .io_in_flow(PE_Array_17_0_io_in_flow),
    .io_in_shift(PE_Array_17_0_io_in_shift),
    .io_out_activate(PE_Array_17_0_io_out_activate),
    .io_out_weight(PE_Array_17_0_io_out_weight),
    .io_out_psum(PE_Array_17_0_io_out_psum)
  );
  basic_PE PE_Array_17_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_1_clock),
    .reset(PE_Array_17_1_reset),
    .io_in_activate(PE_Array_17_1_io_in_activate),
    .io_in_weight(PE_Array_17_1_io_in_weight),
    .io_in_psum(PE_Array_17_1_io_in_psum),
    .io_in_flow(PE_Array_17_1_io_in_flow),
    .io_in_shift(PE_Array_17_1_io_in_shift),
    .io_out_activate(PE_Array_17_1_io_out_activate),
    .io_out_weight(PE_Array_17_1_io_out_weight),
    .io_out_psum(PE_Array_17_1_io_out_psum)
  );
  basic_PE PE_Array_17_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_2_clock),
    .reset(PE_Array_17_2_reset),
    .io_in_activate(PE_Array_17_2_io_in_activate),
    .io_in_weight(PE_Array_17_2_io_in_weight),
    .io_in_psum(PE_Array_17_2_io_in_psum),
    .io_in_flow(PE_Array_17_2_io_in_flow),
    .io_in_shift(PE_Array_17_2_io_in_shift),
    .io_out_activate(PE_Array_17_2_io_out_activate),
    .io_out_weight(PE_Array_17_2_io_out_weight),
    .io_out_psum(PE_Array_17_2_io_out_psum)
  );
  basic_PE PE_Array_17_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_3_clock),
    .reset(PE_Array_17_3_reset),
    .io_in_activate(PE_Array_17_3_io_in_activate),
    .io_in_weight(PE_Array_17_3_io_in_weight),
    .io_in_psum(PE_Array_17_3_io_in_psum),
    .io_in_flow(PE_Array_17_3_io_in_flow),
    .io_in_shift(PE_Array_17_3_io_in_shift),
    .io_out_activate(PE_Array_17_3_io_out_activate),
    .io_out_weight(PE_Array_17_3_io_out_weight),
    .io_out_psum(PE_Array_17_3_io_out_psum)
  );
  basic_PE PE_Array_17_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_4_clock),
    .reset(PE_Array_17_4_reset),
    .io_in_activate(PE_Array_17_4_io_in_activate),
    .io_in_weight(PE_Array_17_4_io_in_weight),
    .io_in_psum(PE_Array_17_4_io_in_psum),
    .io_in_flow(PE_Array_17_4_io_in_flow),
    .io_in_shift(PE_Array_17_4_io_in_shift),
    .io_out_activate(PE_Array_17_4_io_out_activate),
    .io_out_weight(PE_Array_17_4_io_out_weight),
    .io_out_psum(PE_Array_17_4_io_out_psum)
  );
  basic_PE PE_Array_17_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_5_clock),
    .reset(PE_Array_17_5_reset),
    .io_in_activate(PE_Array_17_5_io_in_activate),
    .io_in_weight(PE_Array_17_5_io_in_weight),
    .io_in_psum(PE_Array_17_5_io_in_psum),
    .io_in_flow(PE_Array_17_5_io_in_flow),
    .io_in_shift(PE_Array_17_5_io_in_shift),
    .io_out_activate(PE_Array_17_5_io_out_activate),
    .io_out_weight(PE_Array_17_5_io_out_weight),
    .io_out_psum(PE_Array_17_5_io_out_psum)
  );
  basic_PE PE_Array_17_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_6_clock),
    .reset(PE_Array_17_6_reset),
    .io_in_activate(PE_Array_17_6_io_in_activate),
    .io_in_weight(PE_Array_17_6_io_in_weight),
    .io_in_psum(PE_Array_17_6_io_in_psum),
    .io_in_flow(PE_Array_17_6_io_in_flow),
    .io_in_shift(PE_Array_17_6_io_in_shift),
    .io_out_activate(PE_Array_17_6_io_out_activate),
    .io_out_weight(PE_Array_17_6_io_out_weight),
    .io_out_psum(PE_Array_17_6_io_out_psum)
  );
  basic_PE PE_Array_17_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_7_clock),
    .reset(PE_Array_17_7_reset),
    .io_in_activate(PE_Array_17_7_io_in_activate),
    .io_in_weight(PE_Array_17_7_io_in_weight),
    .io_in_psum(PE_Array_17_7_io_in_psum),
    .io_in_flow(PE_Array_17_7_io_in_flow),
    .io_in_shift(PE_Array_17_7_io_in_shift),
    .io_out_activate(PE_Array_17_7_io_out_activate),
    .io_out_weight(PE_Array_17_7_io_out_weight),
    .io_out_psum(PE_Array_17_7_io_out_psum)
  );
  basic_PE PE_Array_17_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_8_clock),
    .reset(PE_Array_17_8_reset),
    .io_in_activate(PE_Array_17_8_io_in_activate),
    .io_in_weight(PE_Array_17_8_io_in_weight),
    .io_in_psum(PE_Array_17_8_io_in_psum),
    .io_in_flow(PE_Array_17_8_io_in_flow),
    .io_in_shift(PE_Array_17_8_io_in_shift),
    .io_out_activate(PE_Array_17_8_io_out_activate),
    .io_out_weight(PE_Array_17_8_io_out_weight),
    .io_out_psum(PE_Array_17_8_io_out_psum)
  );
  basic_PE PE_Array_17_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_9_clock),
    .reset(PE_Array_17_9_reset),
    .io_in_activate(PE_Array_17_9_io_in_activate),
    .io_in_weight(PE_Array_17_9_io_in_weight),
    .io_in_psum(PE_Array_17_9_io_in_psum),
    .io_in_flow(PE_Array_17_9_io_in_flow),
    .io_in_shift(PE_Array_17_9_io_in_shift),
    .io_out_activate(PE_Array_17_9_io_out_activate),
    .io_out_weight(PE_Array_17_9_io_out_weight),
    .io_out_psum(PE_Array_17_9_io_out_psum)
  );
  basic_PE PE_Array_17_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_10_clock),
    .reset(PE_Array_17_10_reset),
    .io_in_activate(PE_Array_17_10_io_in_activate),
    .io_in_weight(PE_Array_17_10_io_in_weight),
    .io_in_psum(PE_Array_17_10_io_in_psum),
    .io_in_flow(PE_Array_17_10_io_in_flow),
    .io_in_shift(PE_Array_17_10_io_in_shift),
    .io_out_activate(PE_Array_17_10_io_out_activate),
    .io_out_weight(PE_Array_17_10_io_out_weight),
    .io_out_psum(PE_Array_17_10_io_out_psum)
  );
  basic_PE PE_Array_17_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_11_clock),
    .reset(PE_Array_17_11_reset),
    .io_in_activate(PE_Array_17_11_io_in_activate),
    .io_in_weight(PE_Array_17_11_io_in_weight),
    .io_in_psum(PE_Array_17_11_io_in_psum),
    .io_in_flow(PE_Array_17_11_io_in_flow),
    .io_in_shift(PE_Array_17_11_io_in_shift),
    .io_out_activate(PE_Array_17_11_io_out_activate),
    .io_out_weight(PE_Array_17_11_io_out_weight),
    .io_out_psum(PE_Array_17_11_io_out_psum)
  );
  basic_PE PE_Array_17_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_12_clock),
    .reset(PE_Array_17_12_reset),
    .io_in_activate(PE_Array_17_12_io_in_activate),
    .io_in_weight(PE_Array_17_12_io_in_weight),
    .io_in_psum(PE_Array_17_12_io_in_psum),
    .io_in_flow(PE_Array_17_12_io_in_flow),
    .io_in_shift(PE_Array_17_12_io_in_shift),
    .io_out_activate(PE_Array_17_12_io_out_activate),
    .io_out_weight(PE_Array_17_12_io_out_weight),
    .io_out_psum(PE_Array_17_12_io_out_psum)
  );
  basic_PE PE_Array_17_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_13_clock),
    .reset(PE_Array_17_13_reset),
    .io_in_activate(PE_Array_17_13_io_in_activate),
    .io_in_weight(PE_Array_17_13_io_in_weight),
    .io_in_psum(PE_Array_17_13_io_in_psum),
    .io_in_flow(PE_Array_17_13_io_in_flow),
    .io_in_shift(PE_Array_17_13_io_in_shift),
    .io_out_activate(PE_Array_17_13_io_out_activate),
    .io_out_weight(PE_Array_17_13_io_out_weight),
    .io_out_psum(PE_Array_17_13_io_out_psum)
  );
  basic_PE PE_Array_17_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_14_clock),
    .reset(PE_Array_17_14_reset),
    .io_in_activate(PE_Array_17_14_io_in_activate),
    .io_in_weight(PE_Array_17_14_io_in_weight),
    .io_in_psum(PE_Array_17_14_io_in_psum),
    .io_in_flow(PE_Array_17_14_io_in_flow),
    .io_in_shift(PE_Array_17_14_io_in_shift),
    .io_out_activate(PE_Array_17_14_io_out_activate),
    .io_out_weight(PE_Array_17_14_io_out_weight),
    .io_out_psum(PE_Array_17_14_io_out_psum)
  );
  basic_PE PE_Array_17_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_15_clock),
    .reset(PE_Array_17_15_reset),
    .io_in_activate(PE_Array_17_15_io_in_activate),
    .io_in_weight(PE_Array_17_15_io_in_weight),
    .io_in_psum(PE_Array_17_15_io_in_psum),
    .io_in_flow(PE_Array_17_15_io_in_flow),
    .io_in_shift(PE_Array_17_15_io_in_shift),
    .io_out_activate(PE_Array_17_15_io_out_activate),
    .io_out_weight(PE_Array_17_15_io_out_weight),
    .io_out_psum(PE_Array_17_15_io_out_psum)
  );
  basic_PE PE_Array_17_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_16_clock),
    .reset(PE_Array_17_16_reset),
    .io_in_activate(PE_Array_17_16_io_in_activate),
    .io_in_weight(PE_Array_17_16_io_in_weight),
    .io_in_psum(PE_Array_17_16_io_in_psum),
    .io_in_flow(PE_Array_17_16_io_in_flow),
    .io_in_shift(PE_Array_17_16_io_in_shift),
    .io_out_activate(PE_Array_17_16_io_out_activate),
    .io_out_weight(PE_Array_17_16_io_out_weight),
    .io_out_psum(PE_Array_17_16_io_out_psum)
  );
  basic_PE PE_Array_17_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_17_clock),
    .reset(PE_Array_17_17_reset),
    .io_in_activate(PE_Array_17_17_io_in_activate),
    .io_in_weight(PE_Array_17_17_io_in_weight),
    .io_in_psum(PE_Array_17_17_io_in_psum),
    .io_in_flow(PE_Array_17_17_io_in_flow),
    .io_in_shift(PE_Array_17_17_io_in_shift),
    .io_out_activate(PE_Array_17_17_io_out_activate),
    .io_out_weight(PE_Array_17_17_io_out_weight),
    .io_out_psum(PE_Array_17_17_io_out_psum)
  );
  basic_PE PE_Array_17_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_18_clock),
    .reset(PE_Array_17_18_reset),
    .io_in_activate(PE_Array_17_18_io_in_activate),
    .io_in_weight(PE_Array_17_18_io_in_weight),
    .io_in_psum(PE_Array_17_18_io_in_psum),
    .io_in_flow(PE_Array_17_18_io_in_flow),
    .io_in_shift(PE_Array_17_18_io_in_shift),
    .io_out_activate(PE_Array_17_18_io_out_activate),
    .io_out_weight(PE_Array_17_18_io_out_weight),
    .io_out_psum(PE_Array_17_18_io_out_psum)
  );
  basic_PE PE_Array_17_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_19_clock),
    .reset(PE_Array_17_19_reset),
    .io_in_activate(PE_Array_17_19_io_in_activate),
    .io_in_weight(PE_Array_17_19_io_in_weight),
    .io_in_psum(PE_Array_17_19_io_in_psum),
    .io_in_flow(PE_Array_17_19_io_in_flow),
    .io_in_shift(PE_Array_17_19_io_in_shift),
    .io_out_activate(PE_Array_17_19_io_out_activate),
    .io_out_weight(PE_Array_17_19_io_out_weight),
    .io_out_psum(PE_Array_17_19_io_out_psum)
  );
  basic_PE PE_Array_17_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_20_clock),
    .reset(PE_Array_17_20_reset),
    .io_in_activate(PE_Array_17_20_io_in_activate),
    .io_in_weight(PE_Array_17_20_io_in_weight),
    .io_in_psum(PE_Array_17_20_io_in_psum),
    .io_in_flow(PE_Array_17_20_io_in_flow),
    .io_in_shift(PE_Array_17_20_io_in_shift),
    .io_out_activate(PE_Array_17_20_io_out_activate),
    .io_out_weight(PE_Array_17_20_io_out_weight),
    .io_out_psum(PE_Array_17_20_io_out_psum)
  );
  basic_PE PE_Array_17_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_21_clock),
    .reset(PE_Array_17_21_reset),
    .io_in_activate(PE_Array_17_21_io_in_activate),
    .io_in_weight(PE_Array_17_21_io_in_weight),
    .io_in_psum(PE_Array_17_21_io_in_psum),
    .io_in_flow(PE_Array_17_21_io_in_flow),
    .io_in_shift(PE_Array_17_21_io_in_shift),
    .io_out_activate(PE_Array_17_21_io_out_activate),
    .io_out_weight(PE_Array_17_21_io_out_weight),
    .io_out_psum(PE_Array_17_21_io_out_psum)
  );
  basic_PE PE_Array_17_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_22_clock),
    .reset(PE_Array_17_22_reset),
    .io_in_activate(PE_Array_17_22_io_in_activate),
    .io_in_weight(PE_Array_17_22_io_in_weight),
    .io_in_psum(PE_Array_17_22_io_in_psum),
    .io_in_flow(PE_Array_17_22_io_in_flow),
    .io_in_shift(PE_Array_17_22_io_in_shift),
    .io_out_activate(PE_Array_17_22_io_out_activate),
    .io_out_weight(PE_Array_17_22_io_out_weight),
    .io_out_psum(PE_Array_17_22_io_out_psum)
  );
  basic_PE PE_Array_17_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_23_clock),
    .reset(PE_Array_17_23_reset),
    .io_in_activate(PE_Array_17_23_io_in_activate),
    .io_in_weight(PE_Array_17_23_io_in_weight),
    .io_in_psum(PE_Array_17_23_io_in_psum),
    .io_in_flow(PE_Array_17_23_io_in_flow),
    .io_in_shift(PE_Array_17_23_io_in_shift),
    .io_out_activate(PE_Array_17_23_io_out_activate),
    .io_out_weight(PE_Array_17_23_io_out_weight),
    .io_out_psum(PE_Array_17_23_io_out_psum)
  );
  basic_PE PE_Array_17_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_24_clock),
    .reset(PE_Array_17_24_reset),
    .io_in_activate(PE_Array_17_24_io_in_activate),
    .io_in_weight(PE_Array_17_24_io_in_weight),
    .io_in_psum(PE_Array_17_24_io_in_psum),
    .io_in_flow(PE_Array_17_24_io_in_flow),
    .io_in_shift(PE_Array_17_24_io_in_shift),
    .io_out_activate(PE_Array_17_24_io_out_activate),
    .io_out_weight(PE_Array_17_24_io_out_weight),
    .io_out_psum(PE_Array_17_24_io_out_psum)
  );
  basic_PE PE_Array_17_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_25_clock),
    .reset(PE_Array_17_25_reset),
    .io_in_activate(PE_Array_17_25_io_in_activate),
    .io_in_weight(PE_Array_17_25_io_in_weight),
    .io_in_psum(PE_Array_17_25_io_in_psum),
    .io_in_flow(PE_Array_17_25_io_in_flow),
    .io_in_shift(PE_Array_17_25_io_in_shift),
    .io_out_activate(PE_Array_17_25_io_out_activate),
    .io_out_weight(PE_Array_17_25_io_out_weight),
    .io_out_psum(PE_Array_17_25_io_out_psum)
  );
  basic_PE PE_Array_17_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_26_clock),
    .reset(PE_Array_17_26_reset),
    .io_in_activate(PE_Array_17_26_io_in_activate),
    .io_in_weight(PE_Array_17_26_io_in_weight),
    .io_in_psum(PE_Array_17_26_io_in_psum),
    .io_in_flow(PE_Array_17_26_io_in_flow),
    .io_in_shift(PE_Array_17_26_io_in_shift),
    .io_out_activate(PE_Array_17_26_io_out_activate),
    .io_out_weight(PE_Array_17_26_io_out_weight),
    .io_out_psum(PE_Array_17_26_io_out_psum)
  );
  basic_PE PE_Array_17_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_27_clock),
    .reset(PE_Array_17_27_reset),
    .io_in_activate(PE_Array_17_27_io_in_activate),
    .io_in_weight(PE_Array_17_27_io_in_weight),
    .io_in_psum(PE_Array_17_27_io_in_psum),
    .io_in_flow(PE_Array_17_27_io_in_flow),
    .io_in_shift(PE_Array_17_27_io_in_shift),
    .io_out_activate(PE_Array_17_27_io_out_activate),
    .io_out_weight(PE_Array_17_27_io_out_weight),
    .io_out_psum(PE_Array_17_27_io_out_psum)
  );
  basic_PE PE_Array_17_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_28_clock),
    .reset(PE_Array_17_28_reset),
    .io_in_activate(PE_Array_17_28_io_in_activate),
    .io_in_weight(PE_Array_17_28_io_in_weight),
    .io_in_psum(PE_Array_17_28_io_in_psum),
    .io_in_flow(PE_Array_17_28_io_in_flow),
    .io_in_shift(PE_Array_17_28_io_in_shift),
    .io_out_activate(PE_Array_17_28_io_out_activate),
    .io_out_weight(PE_Array_17_28_io_out_weight),
    .io_out_psum(PE_Array_17_28_io_out_psum)
  );
  basic_PE PE_Array_17_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_29_clock),
    .reset(PE_Array_17_29_reset),
    .io_in_activate(PE_Array_17_29_io_in_activate),
    .io_in_weight(PE_Array_17_29_io_in_weight),
    .io_in_psum(PE_Array_17_29_io_in_psum),
    .io_in_flow(PE_Array_17_29_io_in_flow),
    .io_in_shift(PE_Array_17_29_io_in_shift),
    .io_out_activate(PE_Array_17_29_io_out_activate),
    .io_out_weight(PE_Array_17_29_io_out_weight),
    .io_out_psum(PE_Array_17_29_io_out_psum)
  );
  basic_PE PE_Array_17_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_30_clock),
    .reset(PE_Array_17_30_reset),
    .io_in_activate(PE_Array_17_30_io_in_activate),
    .io_in_weight(PE_Array_17_30_io_in_weight),
    .io_in_psum(PE_Array_17_30_io_in_psum),
    .io_in_flow(PE_Array_17_30_io_in_flow),
    .io_in_shift(PE_Array_17_30_io_in_shift),
    .io_out_activate(PE_Array_17_30_io_out_activate),
    .io_out_weight(PE_Array_17_30_io_out_weight),
    .io_out_psum(PE_Array_17_30_io_out_psum)
  );
  basic_PE PE_Array_17_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_17_31_clock),
    .reset(PE_Array_17_31_reset),
    .io_in_activate(PE_Array_17_31_io_in_activate),
    .io_in_weight(PE_Array_17_31_io_in_weight),
    .io_in_psum(PE_Array_17_31_io_in_psum),
    .io_in_flow(PE_Array_17_31_io_in_flow),
    .io_in_shift(PE_Array_17_31_io_in_shift),
    .io_out_activate(PE_Array_17_31_io_out_activate),
    .io_out_weight(PE_Array_17_31_io_out_weight),
    .io_out_psum(PE_Array_17_31_io_out_psum)
  );
  basic_PE PE_Array_18_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_0_clock),
    .reset(PE_Array_18_0_reset),
    .io_in_activate(PE_Array_18_0_io_in_activate),
    .io_in_weight(PE_Array_18_0_io_in_weight),
    .io_in_psum(PE_Array_18_0_io_in_psum),
    .io_in_flow(PE_Array_18_0_io_in_flow),
    .io_in_shift(PE_Array_18_0_io_in_shift),
    .io_out_activate(PE_Array_18_0_io_out_activate),
    .io_out_weight(PE_Array_18_0_io_out_weight),
    .io_out_psum(PE_Array_18_0_io_out_psum)
  );
  basic_PE PE_Array_18_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_1_clock),
    .reset(PE_Array_18_1_reset),
    .io_in_activate(PE_Array_18_1_io_in_activate),
    .io_in_weight(PE_Array_18_1_io_in_weight),
    .io_in_psum(PE_Array_18_1_io_in_psum),
    .io_in_flow(PE_Array_18_1_io_in_flow),
    .io_in_shift(PE_Array_18_1_io_in_shift),
    .io_out_activate(PE_Array_18_1_io_out_activate),
    .io_out_weight(PE_Array_18_1_io_out_weight),
    .io_out_psum(PE_Array_18_1_io_out_psum)
  );
  basic_PE PE_Array_18_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_2_clock),
    .reset(PE_Array_18_2_reset),
    .io_in_activate(PE_Array_18_2_io_in_activate),
    .io_in_weight(PE_Array_18_2_io_in_weight),
    .io_in_psum(PE_Array_18_2_io_in_psum),
    .io_in_flow(PE_Array_18_2_io_in_flow),
    .io_in_shift(PE_Array_18_2_io_in_shift),
    .io_out_activate(PE_Array_18_2_io_out_activate),
    .io_out_weight(PE_Array_18_2_io_out_weight),
    .io_out_psum(PE_Array_18_2_io_out_psum)
  );
  basic_PE PE_Array_18_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_3_clock),
    .reset(PE_Array_18_3_reset),
    .io_in_activate(PE_Array_18_3_io_in_activate),
    .io_in_weight(PE_Array_18_3_io_in_weight),
    .io_in_psum(PE_Array_18_3_io_in_psum),
    .io_in_flow(PE_Array_18_3_io_in_flow),
    .io_in_shift(PE_Array_18_3_io_in_shift),
    .io_out_activate(PE_Array_18_3_io_out_activate),
    .io_out_weight(PE_Array_18_3_io_out_weight),
    .io_out_psum(PE_Array_18_3_io_out_psum)
  );
  basic_PE PE_Array_18_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_4_clock),
    .reset(PE_Array_18_4_reset),
    .io_in_activate(PE_Array_18_4_io_in_activate),
    .io_in_weight(PE_Array_18_4_io_in_weight),
    .io_in_psum(PE_Array_18_4_io_in_psum),
    .io_in_flow(PE_Array_18_4_io_in_flow),
    .io_in_shift(PE_Array_18_4_io_in_shift),
    .io_out_activate(PE_Array_18_4_io_out_activate),
    .io_out_weight(PE_Array_18_4_io_out_weight),
    .io_out_psum(PE_Array_18_4_io_out_psum)
  );
  basic_PE PE_Array_18_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_5_clock),
    .reset(PE_Array_18_5_reset),
    .io_in_activate(PE_Array_18_5_io_in_activate),
    .io_in_weight(PE_Array_18_5_io_in_weight),
    .io_in_psum(PE_Array_18_5_io_in_psum),
    .io_in_flow(PE_Array_18_5_io_in_flow),
    .io_in_shift(PE_Array_18_5_io_in_shift),
    .io_out_activate(PE_Array_18_5_io_out_activate),
    .io_out_weight(PE_Array_18_5_io_out_weight),
    .io_out_psum(PE_Array_18_5_io_out_psum)
  );
  basic_PE PE_Array_18_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_6_clock),
    .reset(PE_Array_18_6_reset),
    .io_in_activate(PE_Array_18_6_io_in_activate),
    .io_in_weight(PE_Array_18_6_io_in_weight),
    .io_in_psum(PE_Array_18_6_io_in_psum),
    .io_in_flow(PE_Array_18_6_io_in_flow),
    .io_in_shift(PE_Array_18_6_io_in_shift),
    .io_out_activate(PE_Array_18_6_io_out_activate),
    .io_out_weight(PE_Array_18_6_io_out_weight),
    .io_out_psum(PE_Array_18_6_io_out_psum)
  );
  basic_PE PE_Array_18_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_7_clock),
    .reset(PE_Array_18_7_reset),
    .io_in_activate(PE_Array_18_7_io_in_activate),
    .io_in_weight(PE_Array_18_7_io_in_weight),
    .io_in_psum(PE_Array_18_7_io_in_psum),
    .io_in_flow(PE_Array_18_7_io_in_flow),
    .io_in_shift(PE_Array_18_7_io_in_shift),
    .io_out_activate(PE_Array_18_7_io_out_activate),
    .io_out_weight(PE_Array_18_7_io_out_weight),
    .io_out_psum(PE_Array_18_7_io_out_psum)
  );
  basic_PE PE_Array_18_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_8_clock),
    .reset(PE_Array_18_8_reset),
    .io_in_activate(PE_Array_18_8_io_in_activate),
    .io_in_weight(PE_Array_18_8_io_in_weight),
    .io_in_psum(PE_Array_18_8_io_in_psum),
    .io_in_flow(PE_Array_18_8_io_in_flow),
    .io_in_shift(PE_Array_18_8_io_in_shift),
    .io_out_activate(PE_Array_18_8_io_out_activate),
    .io_out_weight(PE_Array_18_8_io_out_weight),
    .io_out_psum(PE_Array_18_8_io_out_psum)
  );
  basic_PE PE_Array_18_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_9_clock),
    .reset(PE_Array_18_9_reset),
    .io_in_activate(PE_Array_18_9_io_in_activate),
    .io_in_weight(PE_Array_18_9_io_in_weight),
    .io_in_psum(PE_Array_18_9_io_in_psum),
    .io_in_flow(PE_Array_18_9_io_in_flow),
    .io_in_shift(PE_Array_18_9_io_in_shift),
    .io_out_activate(PE_Array_18_9_io_out_activate),
    .io_out_weight(PE_Array_18_9_io_out_weight),
    .io_out_psum(PE_Array_18_9_io_out_psum)
  );
  basic_PE PE_Array_18_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_10_clock),
    .reset(PE_Array_18_10_reset),
    .io_in_activate(PE_Array_18_10_io_in_activate),
    .io_in_weight(PE_Array_18_10_io_in_weight),
    .io_in_psum(PE_Array_18_10_io_in_psum),
    .io_in_flow(PE_Array_18_10_io_in_flow),
    .io_in_shift(PE_Array_18_10_io_in_shift),
    .io_out_activate(PE_Array_18_10_io_out_activate),
    .io_out_weight(PE_Array_18_10_io_out_weight),
    .io_out_psum(PE_Array_18_10_io_out_psum)
  );
  basic_PE PE_Array_18_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_11_clock),
    .reset(PE_Array_18_11_reset),
    .io_in_activate(PE_Array_18_11_io_in_activate),
    .io_in_weight(PE_Array_18_11_io_in_weight),
    .io_in_psum(PE_Array_18_11_io_in_psum),
    .io_in_flow(PE_Array_18_11_io_in_flow),
    .io_in_shift(PE_Array_18_11_io_in_shift),
    .io_out_activate(PE_Array_18_11_io_out_activate),
    .io_out_weight(PE_Array_18_11_io_out_weight),
    .io_out_psum(PE_Array_18_11_io_out_psum)
  );
  basic_PE PE_Array_18_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_12_clock),
    .reset(PE_Array_18_12_reset),
    .io_in_activate(PE_Array_18_12_io_in_activate),
    .io_in_weight(PE_Array_18_12_io_in_weight),
    .io_in_psum(PE_Array_18_12_io_in_psum),
    .io_in_flow(PE_Array_18_12_io_in_flow),
    .io_in_shift(PE_Array_18_12_io_in_shift),
    .io_out_activate(PE_Array_18_12_io_out_activate),
    .io_out_weight(PE_Array_18_12_io_out_weight),
    .io_out_psum(PE_Array_18_12_io_out_psum)
  );
  basic_PE PE_Array_18_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_13_clock),
    .reset(PE_Array_18_13_reset),
    .io_in_activate(PE_Array_18_13_io_in_activate),
    .io_in_weight(PE_Array_18_13_io_in_weight),
    .io_in_psum(PE_Array_18_13_io_in_psum),
    .io_in_flow(PE_Array_18_13_io_in_flow),
    .io_in_shift(PE_Array_18_13_io_in_shift),
    .io_out_activate(PE_Array_18_13_io_out_activate),
    .io_out_weight(PE_Array_18_13_io_out_weight),
    .io_out_psum(PE_Array_18_13_io_out_psum)
  );
  basic_PE PE_Array_18_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_14_clock),
    .reset(PE_Array_18_14_reset),
    .io_in_activate(PE_Array_18_14_io_in_activate),
    .io_in_weight(PE_Array_18_14_io_in_weight),
    .io_in_psum(PE_Array_18_14_io_in_psum),
    .io_in_flow(PE_Array_18_14_io_in_flow),
    .io_in_shift(PE_Array_18_14_io_in_shift),
    .io_out_activate(PE_Array_18_14_io_out_activate),
    .io_out_weight(PE_Array_18_14_io_out_weight),
    .io_out_psum(PE_Array_18_14_io_out_psum)
  );
  basic_PE PE_Array_18_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_15_clock),
    .reset(PE_Array_18_15_reset),
    .io_in_activate(PE_Array_18_15_io_in_activate),
    .io_in_weight(PE_Array_18_15_io_in_weight),
    .io_in_psum(PE_Array_18_15_io_in_psum),
    .io_in_flow(PE_Array_18_15_io_in_flow),
    .io_in_shift(PE_Array_18_15_io_in_shift),
    .io_out_activate(PE_Array_18_15_io_out_activate),
    .io_out_weight(PE_Array_18_15_io_out_weight),
    .io_out_psum(PE_Array_18_15_io_out_psum)
  );
  basic_PE PE_Array_18_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_16_clock),
    .reset(PE_Array_18_16_reset),
    .io_in_activate(PE_Array_18_16_io_in_activate),
    .io_in_weight(PE_Array_18_16_io_in_weight),
    .io_in_psum(PE_Array_18_16_io_in_psum),
    .io_in_flow(PE_Array_18_16_io_in_flow),
    .io_in_shift(PE_Array_18_16_io_in_shift),
    .io_out_activate(PE_Array_18_16_io_out_activate),
    .io_out_weight(PE_Array_18_16_io_out_weight),
    .io_out_psum(PE_Array_18_16_io_out_psum)
  );
  basic_PE PE_Array_18_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_17_clock),
    .reset(PE_Array_18_17_reset),
    .io_in_activate(PE_Array_18_17_io_in_activate),
    .io_in_weight(PE_Array_18_17_io_in_weight),
    .io_in_psum(PE_Array_18_17_io_in_psum),
    .io_in_flow(PE_Array_18_17_io_in_flow),
    .io_in_shift(PE_Array_18_17_io_in_shift),
    .io_out_activate(PE_Array_18_17_io_out_activate),
    .io_out_weight(PE_Array_18_17_io_out_weight),
    .io_out_psum(PE_Array_18_17_io_out_psum)
  );
  basic_PE PE_Array_18_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_18_clock),
    .reset(PE_Array_18_18_reset),
    .io_in_activate(PE_Array_18_18_io_in_activate),
    .io_in_weight(PE_Array_18_18_io_in_weight),
    .io_in_psum(PE_Array_18_18_io_in_psum),
    .io_in_flow(PE_Array_18_18_io_in_flow),
    .io_in_shift(PE_Array_18_18_io_in_shift),
    .io_out_activate(PE_Array_18_18_io_out_activate),
    .io_out_weight(PE_Array_18_18_io_out_weight),
    .io_out_psum(PE_Array_18_18_io_out_psum)
  );
  basic_PE PE_Array_18_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_19_clock),
    .reset(PE_Array_18_19_reset),
    .io_in_activate(PE_Array_18_19_io_in_activate),
    .io_in_weight(PE_Array_18_19_io_in_weight),
    .io_in_psum(PE_Array_18_19_io_in_psum),
    .io_in_flow(PE_Array_18_19_io_in_flow),
    .io_in_shift(PE_Array_18_19_io_in_shift),
    .io_out_activate(PE_Array_18_19_io_out_activate),
    .io_out_weight(PE_Array_18_19_io_out_weight),
    .io_out_psum(PE_Array_18_19_io_out_psum)
  );
  basic_PE PE_Array_18_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_20_clock),
    .reset(PE_Array_18_20_reset),
    .io_in_activate(PE_Array_18_20_io_in_activate),
    .io_in_weight(PE_Array_18_20_io_in_weight),
    .io_in_psum(PE_Array_18_20_io_in_psum),
    .io_in_flow(PE_Array_18_20_io_in_flow),
    .io_in_shift(PE_Array_18_20_io_in_shift),
    .io_out_activate(PE_Array_18_20_io_out_activate),
    .io_out_weight(PE_Array_18_20_io_out_weight),
    .io_out_psum(PE_Array_18_20_io_out_psum)
  );
  basic_PE PE_Array_18_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_21_clock),
    .reset(PE_Array_18_21_reset),
    .io_in_activate(PE_Array_18_21_io_in_activate),
    .io_in_weight(PE_Array_18_21_io_in_weight),
    .io_in_psum(PE_Array_18_21_io_in_psum),
    .io_in_flow(PE_Array_18_21_io_in_flow),
    .io_in_shift(PE_Array_18_21_io_in_shift),
    .io_out_activate(PE_Array_18_21_io_out_activate),
    .io_out_weight(PE_Array_18_21_io_out_weight),
    .io_out_psum(PE_Array_18_21_io_out_psum)
  );
  basic_PE PE_Array_18_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_22_clock),
    .reset(PE_Array_18_22_reset),
    .io_in_activate(PE_Array_18_22_io_in_activate),
    .io_in_weight(PE_Array_18_22_io_in_weight),
    .io_in_psum(PE_Array_18_22_io_in_psum),
    .io_in_flow(PE_Array_18_22_io_in_flow),
    .io_in_shift(PE_Array_18_22_io_in_shift),
    .io_out_activate(PE_Array_18_22_io_out_activate),
    .io_out_weight(PE_Array_18_22_io_out_weight),
    .io_out_psum(PE_Array_18_22_io_out_psum)
  );
  basic_PE PE_Array_18_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_23_clock),
    .reset(PE_Array_18_23_reset),
    .io_in_activate(PE_Array_18_23_io_in_activate),
    .io_in_weight(PE_Array_18_23_io_in_weight),
    .io_in_psum(PE_Array_18_23_io_in_psum),
    .io_in_flow(PE_Array_18_23_io_in_flow),
    .io_in_shift(PE_Array_18_23_io_in_shift),
    .io_out_activate(PE_Array_18_23_io_out_activate),
    .io_out_weight(PE_Array_18_23_io_out_weight),
    .io_out_psum(PE_Array_18_23_io_out_psum)
  );
  basic_PE PE_Array_18_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_24_clock),
    .reset(PE_Array_18_24_reset),
    .io_in_activate(PE_Array_18_24_io_in_activate),
    .io_in_weight(PE_Array_18_24_io_in_weight),
    .io_in_psum(PE_Array_18_24_io_in_psum),
    .io_in_flow(PE_Array_18_24_io_in_flow),
    .io_in_shift(PE_Array_18_24_io_in_shift),
    .io_out_activate(PE_Array_18_24_io_out_activate),
    .io_out_weight(PE_Array_18_24_io_out_weight),
    .io_out_psum(PE_Array_18_24_io_out_psum)
  );
  basic_PE PE_Array_18_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_25_clock),
    .reset(PE_Array_18_25_reset),
    .io_in_activate(PE_Array_18_25_io_in_activate),
    .io_in_weight(PE_Array_18_25_io_in_weight),
    .io_in_psum(PE_Array_18_25_io_in_psum),
    .io_in_flow(PE_Array_18_25_io_in_flow),
    .io_in_shift(PE_Array_18_25_io_in_shift),
    .io_out_activate(PE_Array_18_25_io_out_activate),
    .io_out_weight(PE_Array_18_25_io_out_weight),
    .io_out_psum(PE_Array_18_25_io_out_psum)
  );
  basic_PE PE_Array_18_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_26_clock),
    .reset(PE_Array_18_26_reset),
    .io_in_activate(PE_Array_18_26_io_in_activate),
    .io_in_weight(PE_Array_18_26_io_in_weight),
    .io_in_psum(PE_Array_18_26_io_in_psum),
    .io_in_flow(PE_Array_18_26_io_in_flow),
    .io_in_shift(PE_Array_18_26_io_in_shift),
    .io_out_activate(PE_Array_18_26_io_out_activate),
    .io_out_weight(PE_Array_18_26_io_out_weight),
    .io_out_psum(PE_Array_18_26_io_out_psum)
  );
  basic_PE PE_Array_18_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_27_clock),
    .reset(PE_Array_18_27_reset),
    .io_in_activate(PE_Array_18_27_io_in_activate),
    .io_in_weight(PE_Array_18_27_io_in_weight),
    .io_in_psum(PE_Array_18_27_io_in_psum),
    .io_in_flow(PE_Array_18_27_io_in_flow),
    .io_in_shift(PE_Array_18_27_io_in_shift),
    .io_out_activate(PE_Array_18_27_io_out_activate),
    .io_out_weight(PE_Array_18_27_io_out_weight),
    .io_out_psum(PE_Array_18_27_io_out_psum)
  );
  basic_PE PE_Array_18_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_28_clock),
    .reset(PE_Array_18_28_reset),
    .io_in_activate(PE_Array_18_28_io_in_activate),
    .io_in_weight(PE_Array_18_28_io_in_weight),
    .io_in_psum(PE_Array_18_28_io_in_psum),
    .io_in_flow(PE_Array_18_28_io_in_flow),
    .io_in_shift(PE_Array_18_28_io_in_shift),
    .io_out_activate(PE_Array_18_28_io_out_activate),
    .io_out_weight(PE_Array_18_28_io_out_weight),
    .io_out_psum(PE_Array_18_28_io_out_psum)
  );
  basic_PE PE_Array_18_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_29_clock),
    .reset(PE_Array_18_29_reset),
    .io_in_activate(PE_Array_18_29_io_in_activate),
    .io_in_weight(PE_Array_18_29_io_in_weight),
    .io_in_psum(PE_Array_18_29_io_in_psum),
    .io_in_flow(PE_Array_18_29_io_in_flow),
    .io_in_shift(PE_Array_18_29_io_in_shift),
    .io_out_activate(PE_Array_18_29_io_out_activate),
    .io_out_weight(PE_Array_18_29_io_out_weight),
    .io_out_psum(PE_Array_18_29_io_out_psum)
  );
  basic_PE PE_Array_18_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_30_clock),
    .reset(PE_Array_18_30_reset),
    .io_in_activate(PE_Array_18_30_io_in_activate),
    .io_in_weight(PE_Array_18_30_io_in_weight),
    .io_in_psum(PE_Array_18_30_io_in_psum),
    .io_in_flow(PE_Array_18_30_io_in_flow),
    .io_in_shift(PE_Array_18_30_io_in_shift),
    .io_out_activate(PE_Array_18_30_io_out_activate),
    .io_out_weight(PE_Array_18_30_io_out_weight),
    .io_out_psum(PE_Array_18_30_io_out_psum)
  );
  basic_PE PE_Array_18_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_18_31_clock),
    .reset(PE_Array_18_31_reset),
    .io_in_activate(PE_Array_18_31_io_in_activate),
    .io_in_weight(PE_Array_18_31_io_in_weight),
    .io_in_psum(PE_Array_18_31_io_in_psum),
    .io_in_flow(PE_Array_18_31_io_in_flow),
    .io_in_shift(PE_Array_18_31_io_in_shift),
    .io_out_activate(PE_Array_18_31_io_out_activate),
    .io_out_weight(PE_Array_18_31_io_out_weight),
    .io_out_psum(PE_Array_18_31_io_out_psum)
  );
  basic_PE PE_Array_19_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_0_clock),
    .reset(PE_Array_19_0_reset),
    .io_in_activate(PE_Array_19_0_io_in_activate),
    .io_in_weight(PE_Array_19_0_io_in_weight),
    .io_in_psum(PE_Array_19_0_io_in_psum),
    .io_in_flow(PE_Array_19_0_io_in_flow),
    .io_in_shift(PE_Array_19_0_io_in_shift),
    .io_out_activate(PE_Array_19_0_io_out_activate),
    .io_out_weight(PE_Array_19_0_io_out_weight),
    .io_out_psum(PE_Array_19_0_io_out_psum)
  );
  basic_PE PE_Array_19_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_1_clock),
    .reset(PE_Array_19_1_reset),
    .io_in_activate(PE_Array_19_1_io_in_activate),
    .io_in_weight(PE_Array_19_1_io_in_weight),
    .io_in_psum(PE_Array_19_1_io_in_psum),
    .io_in_flow(PE_Array_19_1_io_in_flow),
    .io_in_shift(PE_Array_19_1_io_in_shift),
    .io_out_activate(PE_Array_19_1_io_out_activate),
    .io_out_weight(PE_Array_19_1_io_out_weight),
    .io_out_psum(PE_Array_19_1_io_out_psum)
  );
  basic_PE PE_Array_19_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_2_clock),
    .reset(PE_Array_19_2_reset),
    .io_in_activate(PE_Array_19_2_io_in_activate),
    .io_in_weight(PE_Array_19_2_io_in_weight),
    .io_in_psum(PE_Array_19_2_io_in_psum),
    .io_in_flow(PE_Array_19_2_io_in_flow),
    .io_in_shift(PE_Array_19_2_io_in_shift),
    .io_out_activate(PE_Array_19_2_io_out_activate),
    .io_out_weight(PE_Array_19_2_io_out_weight),
    .io_out_psum(PE_Array_19_2_io_out_psum)
  );
  basic_PE PE_Array_19_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_3_clock),
    .reset(PE_Array_19_3_reset),
    .io_in_activate(PE_Array_19_3_io_in_activate),
    .io_in_weight(PE_Array_19_3_io_in_weight),
    .io_in_psum(PE_Array_19_3_io_in_psum),
    .io_in_flow(PE_Array_19_3_io_in_flow),
    .io_in_shift(PE_Array_19_3_io_in_shift),
    .io_out_activate(PE_Array_19_3_io_out_activate),
    .io_out_weight(PE_Array_19_3_io_out_weight),
    .io_out_psum(PE_Array_19_3_io_out_psum)
  );
  basic_PE PE_Array_19_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_4_clock),
    .reset(PE_Array_19_4_reset),
    .io_in_activate(PE_Array_19_4_io_in_activate),
    .io_in_weight(PE_Array_19_4_io_in_weight),
    .io_in_psum(PE_Array_19_4_io_in_psum),
    .io_in_flow(PE_Array_19_4_io_in_flow),
    .io_in_shift(PE_Array_19_4_io_in_shift),
    .io_out_activate(PE_Array_19_4_io_out_activate),
    .io_out_weight(PE_Array_19_4_io_out_weight),
    .io_out_psum(PE_Array_19_4_io_out_psum)
  );
  basic_PE PE_Array_19_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_5_clock),
    .reset(PE_Array_19_5_reset),
    .io_in_activate(PE_Array_19_5_io_in_activate),
    .io_in_weight(PE_Array_19_5_io_in_weight),
    .io_in_psum(PE_Array_19_5_io_in_psum),
    .io_in_flow(PE_Array_19_5_io_in_flow),
    .io_in_shift(PE_Array_19_5_io_in_shift),
    .io_out_activate(PE_Array_19_5_io_out_activate),
    .io_out_weight(PE_Array_19_5_io_out_weight),
    .io_out_psum(PE_Array_19_5_io_out_psum)
  );
  basic_PE PE_Array_19_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_6_clock),
    .reset(PE_Array_19_6_reset),
    .io_in_activate(PE_Array_19_6_io_in_activate),
    .io_in_weight(PE_Array_19_6_io_in_weight),
    .io_in_psum(PE_Array_19_6_io_in_psum),
    .io_in_flow(PE_Array_19_6_io_in_flow),
    .io_in_shift(PE_Array_19_6_io_in_shift),
    .io_out_activate(PE_Array_19_6_io_out_activate),
    .io_out_weight(PE_Array_19_6_io_out_weight),
    .io_out_psum(PE_Array_19_6_io_out_psum)
  );
  basic_PE PE_Array_19_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_7_clock),
    .reset(PE_Array_19_7_reset),
    .io_in_activate(PE_Array_19_7_io_in_activate),
    .io_in_weight(PE_Array_19_7_io_in_weight),
    .io_in_psum(PE_Array_19_7_io_in_psum),
    .io_in_flow(PE_Array_19_7_io_in_flow),
    .io_in_shift(PE_Array_19_7_io_in_shift),
    .io_out_activate(PE_Array_19_7_io_out_activate),
    .io_out_weight(PE_Array_19_7_io_out_weight),
    .io_out_psum(PE_Array_19_7_io_out_psum)
  );
  basic_PE PE_Array_19_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_8_clock),
    .reset(PE_Array_19_8_reset),
    .io_in_activate(PE_Array_19_8_io_in_activate),
    .io_in_weight(PE_Array_19_8_io_in_weight),
    .io_in_psum(PE_Array_19_8_io_in_psum),
    .io_in_flow(PE_Array_19_8_io_in_flow),
    .io_in_shift(PE_Array_19_8_io_in_shift),
    .io_out_activate(PE_Array_19_8_io_out_activate),
    .io_out_weight(PE_Array_19_8_io_out_weight),
    .io_out_psum(PE_Array_19_8_io_out_psum)
  );
  basic_PE PE_Array_19_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_9_clock),
    .reset(PE_Array_19_9_reset),
    .io_in_activate(PE_Array_19_9_io_in_activate),
    .io_in_weight(PE_Array_19_9_io_in_weight),
    .io_in_psum(PE_Array_19_9_io_in_psum),
    .io_in_flow(PE_Array_19_9_io_in_flow),
    .io_in_shift(PE_Array_19_9_io_in_shift),
    .io_out_activate(PE_Array_19_9_io_out_activate),
    .io_out_weight(PE_Array_19_9_io_out_weight),
    .io_out_psum(PE_Array_19_9_io_out_psum)
  );
  basic_PE PE_Array_19_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_10_clock),
    .reset(PE_Array_19_10_reset),
    .io_in_activate(PE_Array_19_10_io_in_activate),
    .io_in_weight(PE_Array_19_10_io_in_weight),
    .io_in_psum(PE_Array_19_10_io_in_psum),
    .io_in_flow(PE_Array_19_10_io_in_flow),
    .io_in_shift(PE_Array_19_10_io_in_shift),
    .io_out_activate(PE_Array_19_10_io_out_activate),
    .io_out_weight(PE_Array_19_10_io_out_weight),
    .io_out_psum(PE_Array_19_10_io_out_psum)
  );
  basic_PE PE_Array_19_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_11_clock),
    .reset(PE_Array_19_11_reset),
    .io_in_activate(PE_Array_19_11_io_in_activate),
    .io_in_weight(PE_Array_19_11_io_in_weight),
    .io_in_psum(PE_Array_19_11_io_in_psum),
    .io_in_flow(PE_Array_19_11_io_in_flow),
    .io_in_shift(PE_Array_19_11_io_in_shift),
    .io_out_activate(PE_Array_19_11_io_out_activate),
    .io_out_weight(PE_Array_19_11_io_out_weight),
    .io_out_psum(PE_Array_19_11_io_out_psum)
  );
  basic_PE PE_Array_19_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_12_clock),
    .reset(PE_Array_19_12_reset),
    .io_in_activate(PE_Array_19_12_io_in_activate),
    .io_in_weight(PE_Array_19_12_io_in_weight),
    .io_in_psum(PE_Array_19_12_io_in_psum),
    .io_in_flow(PE_Array_19_12_io_in_flow),
    .io_in_shift(PE_Array_19_12_io_in_shift),
    .io_out_activate(PE_Array_19_12_io_out_activate),
    .io_out_weight(PE_Array_19_12_io_out_weight),
    .io_out_psum(PE_Array_19_12_io_out_psum)
  );
  basic_PE PE_Array_19_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_13_clock),
    .reset(PE_Array_19_13_reset),
    .io_in_activate(PE_Array_19_13_io_in_activate),
    .io_in_weight(PE_Array_19_13_io_in_weight),
    .io_in_psum(PE_Array_19_13_io_in_psum),
    .io_in_flow(PE_Array_19_13_io_in_flow),
    .io_in_shift(PE_Array_19_13_io_in_shift),
    .io_out_activate(PE_Array_19_13_io_out_activate),
    .io_out_weight(PE_Array_19_13_io_out_weight),
    .io_out_psum(PE_Array_19_13_io_out_psum)
  );
  basic_PE PE_Array_19_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_14_clock),
    .reset(PE_Array_19_14_reset),
    .io_in_activate(PE_Array_19_14_io_in_activate),
    .io_in_weight(PE_Array_19_14_io_in_weight),
    .io_in_psum(PE_Array_19_14_io_in_psum),
    .io_in_flow(PE_Array_19_14_io_in_flow),
    .io_in_shift(PE_Array_19_14_io_in_shift),
    .io_out_activate(PE_Array_19_14_io_out_activate),
    .io_out_weight(PE_Array_19_14_io_out_weight),
    .io_out_psum(PE_Array_19_14_io_out_psum)
  );
  basic_PE PE_Array_19_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_15_clock),
    .reset(PE_Array_19_15_reset),
    .io_in_activate(PE_Array_19_15_io_in_activate),
    .io_in_weight(PE_Array_19_15_io_in_weight),
    .io_in_psum(PE_Array_19_15_io_in_psum),
    .io_in_flow(PE_Array_19_15_io_in_flow),
    .io_in_shift(PE_Array_19_15_io_in_shift),
    .io_out_activate(PE_Array_19_15_io_out_activate),
    .io_out_weight(PE_Array_19_15_io_out_weight),
    .io_out_psum(PE_Array_19_15_io_out_psum)
  );
  basic_PE PE_Array_19_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_16_clock),
    .reset(PE_Array_19_16_reset),
    .io_in_activate(PE_Array_19_16_io_in_activate),
    .io_in_weight(PE_Array_19_16_io_in_weight),
    .io_in_psum(PE_Array_19_16_io_in_psum),
    .io_in_flow(PE_Array_19_16_io_in_flow),
    .io_in_shift(PE_Array_19_16_io_in_shift),
    .io_out_activate(PE_Array_19_16_io_out_activate),
    .io_out_weight(PE_Array_19_16_io_out_weight),
    .io_out_psum(PE_Array_19_16_io_out_psum)
  );
  basic_PE PE_Array_19_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_17_clock),
    .reset(PE_Array_19_17_reset),
    .io_in_activate(PE_Array_19_17_io_in_activate),
    .io_in_weight(PE_Array_19_17_io_in_weight),
    .io_in_psum(PE_Array_19_17_io_in_psum),
    .io_in_flow(PE_Array_19_17_io_in_flow),
    .io_in_shift(PE_Array_19_17_io_in_shift),
    .io_out_activate(PE_Array_19_17_io_out_activate),
    .io_out_weight(PE_Array_19_17_io_out_weight),
    .io_out_psum(PE_Array_19_17_io_out_psum)
  );
  basic_PE PE_Array_19_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_18_clock),
    .reset(PE_Array_19_18_reset),
    .io_in_activate(PE_Array_19_18_io_in_activate),
    .io_in_weight(PE_Array_19_18_io_in_weight),
    .io_in_psum(PE_Array_19_18_io_in_psum),
    .io_in_flow(PE_Array_19_18_io_in_flow),
    .io_in_shift(PE_Array_19_18_io_in_shift),
    .io_out_activate(PE_Array_19_18_io_out_activate),
    .io_out_weight(PE_Array_19_18_io_out_weight),
    .io_out_psum(PE_Array_19_18_io_out_psum)
  );
  basic_PE PE_Array_19_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_19_clock),
    .reset(PE_Array_19_19_reset),
    .io_in_activate(PE_Array_19_19_io_in_activate),
    .io_in_weight(PE_Array_19_19_io_in_weight),
    .io_in_psum(PE_Array_19_19_io_in_psum),
    .io_in_flow(PE_Array_19_19_io_in_flow),
    .io_in_shift(PE_Array_19_19_io_in_shift),
    .io_out_activate(PE_Array_19_19_io_out_activate),
    .io_out_weight(PE_Array_19_19_io_out_weight),
    .io_out_psum(PE_Array_19_19_io_out_psum)
  );
  basic_PE PE_Array_19_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_20_clock),
    .reset(PE_Array_19_20_reset),
    .io_in_activate(PE_Array_19_20_io_in_activate),
    .io_in_weight(PE_Array_19_20_io_in_weight),
    .io_in_psum(PE_Array_19_20_io_in_psum),
    .io_in_flow(PE_Array_19_20_io_in_flow),
    .io_in_shift(PE_Array_19_20_io_in_shift),
    .io_out_activate(PE_Array_19_20_io_out_activate),
    .io_out_weight(PE_Array_19_20_io_out_weight),
    .io_out_psum(PE_Array_19_20_io_out_psum)
  );
  basic_PE PE_Array_19_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_21_clock),
    .reset(PE_Array_19_21_reset),
    .io_in_activate(PE_Array_19_21_io_in_activate),
    .io_in_weight(PE_Array_19_21_io_in_weight),
    .io_in_psum(PE_Array_19_21_io_in_psum),
    .io_in_flow(PE_Array_19_21_io_in_flow),
    .io_in_shift(PE_Array_19_21_io_in_shift),
    .io_out_activate(PE_Array_19_21_io_out_activate),
    .io_out_weight(PE_Array_19_21_io_out_weight),
    .io_out_psum(PE_Array_19_21_io_out_psum)
  );
  basic_PE PE_Array_19_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_22_clock),
    .reset(PE_Array_19_22_reset),
    .io_in_activate(PE_Array_19_22_io_in_activate),
    .io_in_weight(PE_Array_19_22_io_in_weight),
    .io_in_psum(PE_Array_19_22_io_in_psum),
    .io_in_flow(PE_Array_19_22_io_in_flow),
    .io_in_shift(PE_Array_19_22_io_in_shift),
    .io_out_activate(PE_Array_19_22_io_out_activate),
    .io_out_weight(PE_Array_19_22_io_out_weight),
    .io_out_psum(PE_Array_19_22_io_out_psum)
  );
  basic_PE PE_Array_19_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_23_clock),
    .reset(PE_Array_19_23_reset),
    .io_in_activate(PE_Array_19_23_io_in_activate),
    .io_in_weight(PE_Array_19_23_io_in_weight),
    .io_in_psum(PE_Array_19_23_io_in_psum),
    .io_in_flow(PE_Array_19_23_io_in_flow),
    .io_in_shift(PE_Array_19_23_io_in_shift),
    .io_out_activate(PE_Array_19_23_io_out_activate),
    .io_out_weight(PE_Array_19_23_io_out_weight),
    .io_out_psum(PE_Array_19_23_io_out_psum)
  );
  basic_PE PE_Array_19_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_24_clock),
    .reset(PE_Array_19_24_reset),
    .io_in_activate(PE_Array_19_24_io_in_activate),
    .io_in_weight(PE_Array_19_24_io_in_weight),
    .io_in_psum(PE_Array_19_24_io_in_psum),
    .io_in_flow(PE_Array_19_24_io_in_flow),
    .io_in_shift(PE_Array_19_24_io_in_shift),
    .io_out_activate(PE_Array_19_24_io_out_activate),
    .io_out_weight(PE_Array_19_24_io_out_weight),
    .io_out_psum(PE_Array_19_24_io_out_psum)
  );
  basic_PE PE_Array_19_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_25_clock),
    .reset(PE_Array_19_25_reset),
    .io_in_activate(PE_Array_19_25_io_in_activate),
    .io_in_weight(PE_Array_19_25_io_in_weight),
    .io_in_psum(PE_Array_19_25_io_in_psum),
    .io_in_flow(PE_Array_19_25_io_in_flow),
    .io_in_shift(PE_Array_19_25_io_in_shift),
    .io_out_activate(PE_Array_19_25_io_out_activate),
    .io_out_weight(PE_Array_19_25_io_out_weight),
    .io_out_psum(PE_Array_19_25_io_out_psum)
  );
  basic_PE PE_Array_19_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_26_clock),
    .reset(PE_Array_19_26_reset),
    .io_in_activate(PE_Array_19_26_io_in_activate),
    .io_in_weight(PE_Array_19_26_io_in_weight),
    .io_in_psum(PE_Array_19_26_io_in_psum),
    .io_in_flow(PE_Array_19_26_io_in_flow),
    .io_in_shift(PE_Array_19_26_io_in_shift),
    .io_out_activate(PE_Array_19_26_io_out_activate),
    .io_out_weight(PE_Array_19_26_io_out_weight),
    .io_out_psum(PE_Array_19_26_io_out_psum)
  );
  basic_PE PE_Array_19_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_27_clock),
    .reset(PE_Array_19_27_reset),
    .io_in_activate(PE_Array_19_27_io_in_activate),
    .io_in_weight(PE_Array_19_27_io_in_weight),
    .io_in_psum(PE_Array_19_27_io_in_psum),
    .io_in_flow(PE_Array_19_27_io_in_flow),
    .io_in_shift(PE_Array_19_27_io_in_shift),
    .io_out_activate(PE_Array_19_27_io_out_activate),
    .io_out_weight(PE_Array_19_27_io_out_weight),
    .io_out_psum(PE_Array_19_27_io_out_psum)
  );
  basic_PE PE_Array_19_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_28_clock),
    .reset(PE_Array_19_28_reset),
    .io_in_activate(PE_Array_19_28_io_in_activate),
    .io_in_weight(PE_Array_19_28_io_in_weight),
    .io_in_psum(PE_Array_19_28_io_in_psum),
    .io_in_flow(PE_Array_19_28_io_in_flow),
    .io_in_shift(PE_Array_19_28_io_in_shift),
    .io_out_activate(PE_Array_19_28_io_out_activate),
    .io_out_weight(PE_Array_19_28_io_out_weight),
    .io_out_psum(PE_Array_19_28_io_out_psum)
  );
  basic_PE PE_Array_19_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_29_clock),
    .reset(PE_Array_19_29_reset),
    .io_in_activate(PE_Array_19_29_io_in_activate),
    .io_in_weight(PE_Array_19_29_io_in_weight),
    .io_in_psum(PE_Array_19_29_io_in_psum),
    .io_in_flow(PE_Array_19_29_io_in_flow),
    .io_in_shift(PE_Array_19_29_io_in_shift),
    .io_out_activate(PE_Array_19_29_io_out_activate),
    .io_out_weight(PE_Array_19_29_io_out_weight),
    .io_out_psum(PE_Array_19_29_io_out_psum)
  );
  basic_PE PE_Array_19_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_30_clock),
    .reset(PE_Array_19_30_reset),
    .io_in_activate(PE_Array_19_30_io_in_activate),
    .io_in_weight(PE_Array_19_30_io_in_weight),
    .io_in_psum(PE_Array_19_30_io_in_psum),
    .io_in_flow(PE_Array_19_30_io_in_flow),
    .io_in_shift(PE_Array_19_30_io_in_shift),
    .io_out_activate(PE_Array_19_30_io_out_activate),
    .io_out_weight(PE_Array_19_30_io_out_weight),
    .io_out_psum(PE_Array_19_30_io_out_psum)
  );
  basic_PE PE_Array_19_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_19_31_clock),
    .reset(PE_Array_19_31_reset),
    .io_in_activate(PE_Array_19_31_io_in_activate),
    .io_in_weight(PE_Array_19_31_io_in_weight),
    .io_in_psum(PE_Array_19_31_io_in_psum),
    .io_in_flow(PE_Array_19_31_io_in_flow),
    .io_in_shift(PE_Array_19_31_io_in_shift),
    .io_out_activate(PE_Array_19_31_io_out_activate),
    .io_out_weight(PE_Array_19_31_io_out_weight),
    .io_out_psum(PE_Array_19_31_io_out_psum)
  );
  basic_PE PE_Array_20_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_0_clock),
    .reset(PE_Array_20_0_reset),
    .io_in_activate(PE_Array_20_0_io_in_activate),
    .io_in_weight(PE_Array_20_0_io_in_weight),
    .io_in_psum(PE_Array_20_0_io_in_psum),
    .io_in_flow(PE_Array_20_0_io_in_flow),
    .io_in_shift(PE_Array_20_0_io_in_shift),
    .io_out_activate(PE_Array_20_0_io_out_activate),
    .io_out_weight(PE_Array_20_0_io_out_weight),
    .io_out_psum(PE_Array_20_0_io_out_psum)
  );
  basic_PE PE_Array_20_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_1_clock),
    .reset(PE_Array_20_1_reset),
    .io_in_activate(PE_Array_20_1_io_in_activate),
    .io_in_weight(PE_Array_20_1_io_in_weight),
    .io_in_psum(PE_Array_20_1_io_in_psum),
    .io_in_flow(PE_Array_20_1_io_in_flow),
    .io_in_shift(PE_Array_20_1_io_in_shift),
    .io_out_activate(PE_Array_20_1_io_out_activate),
    .io_out_weight(PE_Array_20_1_io_out_weight),
    .io_out_psum(PE_Array_20_1_io_out_psum)
  );
  basic_PE PE_Array_20_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_2_clock),
    .reset(PE_Array_20_2_reset),
    .io_in_activate(PE_Array_20_2_io_in_activate),
    .io_in_weight(PE_Array_20_2_io_in_weight),
    .io_in_psum(PE_Array_20_2_io_in_psum),
    .io_in_flow(PE_Array_20_2_io_in_flow),
    .io_in_shift(PE_Array_20_2_io_in_shift),
    .io_out_activate(PE_Array_20_2_io_out_activate),
    .io_out_weight(PE_Array_20_2_io_out_weight),
    .io_out_psum(PE_Array_20_2_io_out_psum)
  );
  basic_PE PE_Array_20_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_3_clock),
    .reset(PE_Array_20_3_reset),
    .io_in_activate(PE_Array_20_3_io_in_activate),
    .io_in_weight(PE_Array_20_3_io_in_weight),
    .io_in_psum(PE_Array_20_3_io_in_psum),
    .io_in_flow(PE_Array_20_3_io_in_flow),
    .io_in_shift(PE_Array_20_3_io_in_shift),
    .io_out_activate(PE_Array_20_3_io_out_activate),
    .io_out_weight(PE_Array_20_3_io_out_weight),
    .io_out_psum(PE_Array_20_3_io_out_psum)
  );
  basic_PE PE_Array_20_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_4_clock),
    .reset(PE_Array_20_4_reset),
    .io_in_activate(PE_Array_20_4_io_in_activate),
    .io_in_weight(PE_Array_20_4_io_in_weight),
    .io_in_psum(PE_Array_20_4_io_in_psum),
    .io_in_flow(PE_Array_20_4_io_in_flow),
    .io_in_shift(PE_Array_20_4_io_in_shift),
    .io_out_activate(PE_Array_20_4_io_out_activate),
    .io_out_weight(PE_Array_20_4_io_out_weight),
    .io_out_psum(PE_Array_20_4_io_out_psum)
  );
  basic_PE PE_Array_20_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_5_clock),
    .reset(PE_Array_20_5_reset),
    .io_in_activate(PE_Array_20_5_io_in_activate),
    .io_in_weight(PE_Array_20_5_io_in_weight),
    .io_in_psum(PE_Array_20_5_io_in_psum),
    .io_in_flow(PE_Array_20_5_io_in_flow),
    .io_in_shift(PE_Array_20_5_io_in_shift),
    .io_out_activate(PE_Array_20_5_io_out_activate),
    .io_out_weight(PE_Array_20_5_io_out_weight),
    .io_out_psum(PE_Array_20_5_io_out_psum)
  );
  basic_PE PE_Array_20_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_6_clock),
    .reset(PE_Array_20_6_reset),
    .io_in_activate(PE_Array_20_6_io_in_activate),
    .io_in_weight(PE_Array_20_6_io_in_weight),
    .io_in_psum(PE_Array_20_6_io_in_psum),
    .io_in_flow(PE_Array_20_6_io_in_flow),
    .io_in_shift(PE_Array_20_6_io_in_shift),
    .io_out_activate(PE_Array_20_6_io_out_activate),
    .io_out_weight(PE_Array_20_6_io_out_weight),
    .io_out_psum(PE_Array_20_6_io_out_psum)
  );
  basic_PE PE_Array_20_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_7_clock),
    .reset(PE_Array_20_7_reset),
    .io_in_activate(PE_Array_20_7_io_in_activate),
    .io_in_weight(PE_Array_20_7_io_in_weight),
    .io_in_psum(PE_Array_20_7_io_in_psum),
    .io_in_flow(PE_Array_20_7_io_in_flow),
    .io_in_shift(PE_Array_20_7_io_in_shift),
    .io_out_activate(PE_Array_20_7_io_out_activate),
    .io_out_weight(PE_Array_20_7_io_out_weight),
    .io_out_psum(PE_Array_20_7_io_out_psum)
  );
  basic_PE PE_Array_20_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_8_clock),
    .reset(PE_Array_20_8_reset),
    .io_in_activate(PE_Array_20_8_io_in_activate),
    .io_in_weight(PE_Array_20_8_io_in_weight),
    .io_in_psum(PE_Array_20_8_io_in_psum),
    .io_in_flow(PE_Array_20_8_io_in_flow),
    .io_in_shift(PE_Array_20_8_io_in_shift),
    .io_out_activate(PE_Array_20_8_io_out_activate),
    .io_out_weight(PE_Array_20_8_io_out_weight),
    .io_out_psum(PE_Array_20_8_io_out_psum)
  );
  basic_PE PE_Array_20_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_9_clock),
    .reset(PE_Array_20_9_reset),
    .io_in_activate(PE_Array_20_9_io_in_activate),
    .io_in_weight(PE_Array_20_9_io_in_weight),
    .io_in_psum(PE_Array_20_9_io_in_psum),
    .io_in_flow(PE_Array_20_9_io_in_flow),
    .io_in_shift(PE_Array_20_9_io_in_shift),
    .io_out_activate(PE_Array_20_9_io_out_activate),
    .io_out_weight(PE_Array_20_9_io_out_weight),
    .io_out_psum(PE_Array_20_9_io_out_psum)
  );
  basic_PE PE_Array_20_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_10_clock),
    .reset(PE_Array_20_10_reset),
    .io_in_activate(PE_Array_20_10_io_in_activate),
    .io_in_weight(PE_Array_20_10_io_in_weight),
    .io_in_psum(PE_Array_20_10_io_in_psum),
    .io_in_flow(PE_Array_20_10_io_in_flow),
    .io_in_shift(PE_Array_20_10_io_in_shift),
    .io_out_activate(PE_Array_20_10_io_out_activate),
    .io_out_weight(PE_Array_20_10_io_out_weight),
    .io_out_psum(PE_Array_20_10_io_out_psum)
  );
  basic_PE PE_Array_20_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_11_clock),
    .reset(PE_Array_20_11_reset),
    .io_in_activate(PE_Array_20_11_io_in_activate),
    .io_in_weight(PE_Array_20_11_io_in_weight),
    .io_in_psum(PE_Array_20_11_io_in_psum),
    .io_in_flow(PE_Array_20_11_io_in_flow),
    .io_in_shift(PE_Array_20_11_io_in_shift),
    .io_out_activate(PE_Array_20_11_io_out_activate),
    .io_out_weight(PE_Array_20_11_io_out_weight),
    .io_out_psum(PE_Array_20_11_io_out_psum)
  );
  basic_PE PE_Array_20_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_12_clock),
    .reset(PE_Array_20_12_reset),
    .io_in_activate(PE_Array_20_12_io_in_activate),
    .io_in_weight(PE_Array_20_12_io_in_weight),
    .io_in_psum(PE_Array_20_12_io_in_psum),
    .io_in_flow(PE_Array_20_12_io_in_flow),
    .io_in_shift(PE_Array_20_12_io_in_shift),
    .io_out_activate(PE_Array_20_12_io_out_activate),
    .io_out_weight(PE_Array_20_12_io_out_weight),
    .io_out_psum(PE_Array_20_12_io_out_psum)
  );
  basic_PE PE_Array_20_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_13_clock),
    .reset(PE_Array_20_13_reset),
    .io_in_activate(PE_Array_20_13_io_in_activate),
    .io_in_weight(PE_Array_20_13_io_in_weight),
    .io_in_psum(PE_Array_20_13_io_in_psum),
    .io_in_flow(PE_Array_20_13_io_in_flow),
    .io_in_shift(PE_Array_20_13_io_in_shift),
    .io_out_activate(PE_Array_20_13_io_out_activate),
    .io_out_weight(PE_Array_20_13_io_out_weight),
    .io_out_psum(PE_Array_20_13_io_out_psum)
  );
  basic_PE PE_Array_20_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_14_clock),
    .reset(PE_Array_20_14_reset),
    .io_in_activate(PE_Array_20_14_io_in_activate),
    .io_in_weight(PE_Array_20_14_io_in_weight),
    .io_in_psum(PE_Array_20_14_io_in_psum),
    .io_in_flow(PE_Array_20_14_io_in_flow),
    .io_in_shift(PE_Array_20_14_io_in_shift),
    .io_out_activate(PE_Array_20_14_io_out_activate),
    .io_out_weight(PE_Array_20_14_io_out_weight),
    .io_out_psum(PE_Array_20_14_io_out_psum)
  );
  basic_PE PE_Array_20_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_15_clock),
    .reset(PE_Array_20_15_reset),
    .io_in_activate(PE_Array_20_15_io_in_activate),
    .io_in_weight(PE_Array_20_15_io_in_weight),
    .io_in_psum(PE_Array_20_15_io_in_psum),
    .io_in_flow(PE_Array_20_15_io_in_flow),
    .io_in_shift(PE_Array_20_15_io_in_shift),
    .io_out_activate(PE_Array_20_15_io_out_activate),
    .io_out_weight(PE_Array_20_15_io_out_weight),
    .io_out_psum(PE_Array_20_15_io_out_psum)
  );
  basic_PE PE_Array_20_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_16_clock),
    .reset(PE_Array_20_16_reset),
    .io_in_activate(PE_Array_20_16_io_in_activate),
    .io_in_weight(PE_Array_20_16_io_in_weight),
    .io_in_psum(PE_Array_20_16_io_in_psum),
    .io_in_flow(PE_Array_20_16_io_in_flow),
    .io_in_shift(PE_Array_20_16_io_in_shift),
    .io_out_activate(PE_Array_20_16_io_out_activate),
    .io_out_weight(PE_Array_20_16_io_out_weight),
    .io_out_psum(PE_Array_20_16_io_out_psum)
  );
  basic_PE PE_Array_20_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_17_clock),
    .reset(PE_Array_20_17_reset),
    .io_in_activate(PE_Array_20_17_io_in_activate),
    .io_in_weight(PE_Array_20_17_io_in_weight),
    .io_in_psum(PE_Array_20_17_io_in_psum),
    .io_in_flow(PE_Array_20_17_io_in_flow),
    .io_in_shift(PE_Array_20_17_io_in_shift),
    .io_out_activate(PE_Array_20_17_io_out_activate),
    .io_out_weight(PE_Array_20_17_io_out_weight),
    .io_out_psum(PE_Array_20_17_io_out_psum)
  );
  basic_PE PE_Array_20_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_18_clock),
    .reset(PE_Array_20_18_reset),
    .io_in_activate(PE_Array_20_18_io_in_activate),
    .io_in_weight(PE_Array_20_18_io_in_weight),
    .io_in_psum(PE_Array_20_18_io_in_psum),
    .io_in_flow(PE_Array_20_18_io_in_flow),
    .io_in_shift(PE_Array_20_18_io_in_shift),
    .io_out_activate(PE_Array_20_18_io_out_activate),
    .io_out_weight(PE_Array_20_18_io_out_weight),
    .io_out_psum(PE_Array_20_18_io_out_psum)
  );
  basic_PE PE_Array_20_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_19_clock),
    .reset(PE_Array_20_19_reset),
    .io_in_activate(PE_Array_20_19_io_in_activate),
    .io_in_weight(PE_Array_20_19_io_in_weight),
    .io_in_psum(PE_Array_20_19_io_in_psum),
    .io_in_flow(PE_Array_20_19_io_in_flow),
    .io_in_shift(PE_Array_20_19_io_in_shift),
    .io_out_activate(PE_Array_20_19_io_out_activate),
    .io_out_weight(PE_Array_20_19_io_out_weight),
    .io_out_psum(PE_Array_20_19_io_out_psum)
  );
  basic_PE PE_Array_20_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_20_clock),
    .reset(PE_Array_20_20_reset),
    .io_in_activate(PE_Array_20_20_io_in_activate),
    .io_in_weight(PE_Array_20_20_io_in_weight),
    .io_in_psum(PE_Array_20_20_io_in_psum),
    .io_in_flow(PE_Array_20_20_io_in_flow),
    .io_in_shift(PE_Array_20_20_io_in_shift),
    .io_out_activate(PE_Array_20_20_io_out_activate),
    .io_out_weight(PE_Array_20_20_io_out_weight),
    .io_out_psum(PE_Array_20_20_io_out_psum)
  );
  basic_PE PE_Array_20_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_21_clock),
    .reset(PE_Array_20_21_reset),
    .io_in_activate(PE_Array_20_21_io_in_activate),
    .io_in_weight(PE_Array_20_21_io_in_weight),
    .io_in_psum(PE_Array_20_21_io_in_psum),
    .io_in_flow(PE_Array_20_21_io_in_flow),
    .io_in_shift(PE_Array_20_21_io_in_shift),
    .io_out_activate(PE_Array_20_21_io_out_activate),
    .io_out_weight(PE_Array_20_21_io_out_weight),
    .io_out_psum(PE_Array_20_21_io_out_psum)
  );
  basic_PE PE_Array_20_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_22_clock),
    .reset(PE_Array_20_22_reset),
    .io_in_activate(PE_Array_20_22_io_in_activate),
    .io_in_weight(PE_Array_20_22_io_in_weight),
    .io_in_psum(PE_Array_20_22_io_in_psum),
    .io_in_flow(PE_Array_20_22_io_in_flow),
    .io_in_shift(PE_Array_20_22_io_in_shift),
    .io_out_activate(PE_Array_20_22_io_out_activate),
    .io_out_weight(PE_Array_20_22_io_out_weight),
    .io_out_psum(PE_Array_20_22_io_out_psum)
  );
  basic_PE PE_Array_20_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_23_clock),
    .reset(PE_Array_20_23_reset),
    .io_in_activate(PE_Array_20_23_io_in_activate),
    .io_in_weight(PE_Array_20_23_io_in_weight),
    .io_in_psum(PE_Array_20_23_io_in_psum),
    .io_in_flow(PE_Array_20_23_io_in_flow),
    .io_in_shift(PE_Array_20_23_io_in_shift),
    .io_out_activate(PE_Array_20_23_io_out_activate),
    .io_out_weight(PE_Array_20_23_io_out_weight),
    .io_out_psum(PE_Array_20_23_io_out_psum)
  );
  basic_PE PE_Array_20_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_24_clock),
    .reset(PE_Array_20_24_reset),
    .io_in_activate(PE_Array_20_24_io_in_activate),
    .io_in_weight(PE_Array_20_24_io_in_weight),
    .io_in_psum(PE_Array_20_24_io_in_psum),
    .io_in_flow(PE_Array_20_24_io_in_flow),
    .io_in_shift(PE_Array_20_24_io_in_shift),
    .io_out_activate(PE_Array_20_24_io_out_activate),
    .io_out_weight(PE_Array_20_24_io_out_weight),
    .io_out_psum(PE_Array_20_24_io_out_psum)
  );
  basic_PE PE_Array_20_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_25_clock),
    .reset(PE_Array_20_25_reset),
    .io_in_activate(PE_Array_20_25_io_in_activate),
    .io_in_weight(PE_Array_20_25_io_in_weight),
    .io_in_psum(PE_Array_20_25_io_in_psum),
    .io_in_flow(PE_Array_20_25_io_in_flow),
    .io_in_shift(PE_Array_20_25_io_in_shift),
    .io_out_activate(PE_Array_20_25_io_out_activate),
    .io_out_weight(PE_Array_20_25_io_out_weight),
    .io_out_psum(PE_Array_20_25_io_out_psum)
  );
  basic_PE PE_Array_20_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_26_clock),
    .reset(PE_Array_20_26_reset),
    .io_in_activate(PE_Array_20_26_io_in_activate),
    .io_in_weight(PE_Array_20_26_io_in_weight),
    .io_in_psum(PE_Array_20_26_io_in_psum),
    .io_in_flow(PE_Array_20_26_io_in_flow),
    .io_in_shift(PE_Array_20_26_io_in_shift),
    .io_out_activate(PE_Array_20_26_io_out_activate),
    .io_out_weight(PE_Array_20_26_io_out_weight),
    .io_out_psum(PE_Array_20_26_io_out_psum)
  );
  basic_PE PE_Array_20_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_27_clock),
    .reset(PE_Array_20_27_reset),
    .io_in_activate(PE_Array_20_27_io_in_activate),
    .io_in_weight(PE_Array_20_27_io_in_weight),
    .io_in_psum(PE_Array_20_27_io_in_psum),
    .io_in_flow(PE_Array_20_27_io_in_flow),
    .io_in_shift(PE_Array_20_27_io_in_shift),
    .io_out_activate(PE_Array_20_27_io_out_activate),
    .io_out_weight(PE_Array_20_27_io_out_weight),
    .io_out_psum(PE_Array_20_27_io_out_psum)
  );
  basic_PE PE_Array_20_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_28_clock),
    .reset(PE_Array_20_28_reset),
    .io_in_activate(PE_Array_20_28_io_in_activate),
    .io_in_weight(PE_Array_20_28_io_in_weight),
    .io_in_psum(PE_Array_20_28_io_in_psum),
    .io_in_flow(PE_Array_20_28_io_in_flow),
    .io_in_shift(PE_Array_20_28_io_in_shift),
    .io_out_activate(PE_Array_20_28_io_out_activate),
    .io_out_weight(PE_Array_20_28_io_out_weight),
    .io_out_psum(PE_Array_20_28_io_out_psum)
  );
  basic_PE PE_Array_20_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_29_clock),
    .reset(PE_Array_20_29_reset),
    .io_in_activate(PE_Array_20_29_io_in_activate),
    .io_in_weight(PE_Array_20_29_io_in_weight),
    .io_in_psum(PE_Array_20_29_io_in_psum),
    .io_in_flow(PE_Array_20_29_io_in_flow),
    .io_in_shift(PE_Array_20_29_io_in_shift),
    .io_out_activate(PE_Array_20_29_io_out_activate),
    .io_out_weight(PE_Array_20_29_io_out_weight),
    .io_out_psum(PE_Array_20_29_io_out_psum)
  );
  basic_PE PE_Array_20_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_30_clock),
    .reset(PE_Array_20_30_reset),
    .io_in_activate(PE_Array_20_30_io_in_activate),
    .io_in_weight(PE_Array_20_30_io_in_weight),
    .io_in_psum(PE_Array_20_30_io_in_psum),
    .io_in_flow(PE_Array_20_30_io_in_flow),
    .io_in_shift(PE_Array_20_30_io_in_shift),
    .io_out_activate(PE_Array_20_30_io_out_activate),
    .io_out_weight(PE_Array_20_30_io_out_weight),
    .io_out_psum(PE_Array_20_30_io_out_psum)
  );
  basic_PE PE_Array_20_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_20_31_clock),
    .reset(PE_Array_20_31_reset),
    .io_in_activate(PE_Array_20_31_io_in_activate),
    .io_in_weight(PE_Array_20_31_io_in_weight),
    .io_in_psum(PE_Array_20_31_io_in_psum),
    .io_in_flow(PE_Array_20_31_io_in_flow),
    .io_in_shift(PE_Array_20_31_io_in_shift),
    .io_out_activate(PE_Array_20_31_io_out_activate),
    .io_out_weight(PE_Array_20_31_io_out_weight),
    .io_out_psum(PE_Array_20_31_io_out_psum)
  );
  basic_PE PE_Array_21_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_0_clock),
    .reset(PE_Array_21_0_reset),
    .io_in_activate(PE_Array_21_0_io_in_activate),
    .io_in_weight(PE_Array_21_0_io_in_weight),
    .io_in_psum(PE_Array_21_0_io_in_psum),
    .io_in_flow(PE_Array_21_0_io_in_flow),
    .io_in_shift(PE_Array_21_0_io_in_shift),
    .io_out_activate(PE_Array_21_0_io_out_activate),
    .io_out_weight(PE_Array_21_0_io_out_weight),
    .io_out_psum(PE_Array_21_0_io_out_psum)
  );
  basic_PE PE_Array_21_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_1_clock),
    .reset(PE_Array_21_1_reset),
    .io_in_activate(PE_Array_21_1_io_in_activate),
    .io_in_weight(PE_Array_21_1_io_in_weight),
    .io_in_psum(PE_Array_21_1_io_in_psum),
    .io_in_flow(PE_Array_21_1_io_in_flow),
    .io_in_shift(PE_Array_21_1_io_in_shift),
    .io_out_activate(PE_Array_21_1_io_out_activate),
    .io_out_weight(PE_Array_21_1_io_out_weight),
    .io_out_psum(PE_Array_21_1_io_out_psum)
  );
  basic_PE PE_Array_21_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_2_clock),
    .reset(PE_Array_21_2_reset),
    .io_in_activate(PE_Array_21_2_io_in_activate),
    .io_in_weight(PE_Array_21_2_io_in_weight),
    .io_in_psum(PE_Array_21_2_io_in_psum),
    .io_in_flow(PE_Array_21_2_io_in_flow),
    .io_in_shift(PE_Array_21_2_io_in_shift),
    .io_out_activate(PE_Array_21_2_io_out_activate),
    .io_out_weight(PE_Array_21_2_io_out_weight),
    .io_out_psum(PE_Array_21_2_io_out_psum)
  );
  basic_PE PE_Array_21_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_3_clock),
    .reset(PE_Array_21_3_reset),
    .io_in_activate(PE_Array_21_3_io_in_activate),
    .io_in_weight(PE_Array_21_3_io_in_weight),
    .io_in_psum(PE_Array_21_3_io_in_psum),
    .io_in_flow(PE_Array_21_3_io_in_flow),
    .io_in_shift(PE_Array_21_3_io_in_shift),
    .io_out_activate(PE_Array_21_3_io_out_activate),
    .io_out_weight(PE_Array_21_3_io_out_weight),
    .io_out_psum(PE_Array_21_3_io_out_psum)
  );
  basic_PE PE_Array_21_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_4_clock),
    .reset(PE_Array_21_4_reset),
    .io_in_activate(PE_Array_21_4_io_in_activate),
    .io_in_weight(PE_Array_21_4_io_in_weight),
    .io_in_psum(PE_Array_21_4_io_in_psum),
    .io_in_flow(PE_Array_21_4_io_in_flow),
    .io_in_shift(PE_Array_21_4_io_in_shift),
    .io_out_activate(PE_Array_21_4_io_out_activate),
    .io_out_weight(PE_Array_21_4_io_out_weight),
    .io_out_psum(PE_Array_21_4_io_out_psum)
  );
  basic_PE PE_Array_21_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_5_clock),
    .reset(PE_Array_21_5_reset),
    .io_in_activate(PE_Array_21_5_io_in_activate),
    .io_in_weight(PE_Array_21_5_io_in_weight),
    .io_in_psum(PE_Array_21_5_io_in_psum),
    .io_in_flow(PE_Array_21_5_io_in_flow),
    .io_in_shift(PE_Array_21_5_io_in_shift),
    .io_out_activate(PE_Array_21_5_io_out_activate),
    .io_out_weight(PE_Array_21_5_io_out_weight),
    .io_out_psum(PE_Array_21_5_io_out_psum)
  );
  basic_PE PE_Array_21_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_6_clock),
    .reset(PE_Array_21_6_reset),
    .io_in_activate(PE_Array_21_6_io_in_activate),
    .io_in_weight(PE_Array_21_6_io_in_weight),
    .io_in_psum(PE_Array_21_6_io_in_psum),
    .io_in_flow(PE_Array_21_6_io_in_flow),
    .io_in_shift(PE_Array_21_6_io_in_shift),
    .io_out_activate(PE_Array_21_6_io_out_activate),
    .io_out_weight(PE_Array_21_6_io_out_weight),
    .io_out_psum(PE_Array_21_6_io_out_psum)
  );
  basic_PE PE_Array_21_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_7_clock),
    .reset(PE_Array_21_7_reset),
    .io_in_activate(PE_Array_21_7_io_in_activate),
    .io_in_weight(PE_Array_21_7_io_in_weight),
    .io_in_psum(PE_Array_21_7_io_in_psum),
    .io_in_flow(PE_Array_21_7_io_in_flow),
    .io_in_shift(PE_Array_21_7_io_in_shift),
    .io_out_activate(PE_Array_21_7_io_out_activate),
    .io_out_weight(PE_Array_21_7_io_out_weight),
    .io_out_psum(PE_Array_21_7_io_out_psum)
  );
  basic_PE PE_Array_21_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_8_clock),
    .reset(PE_Array_21_8_reset),
    .io_in_activate(PE_Array_21_8_io_in_activate),
    .io_in_weight(PE_Array_21_8_io_in_weight),
    .io_in_psum(PE_Array_21_8_io_in_psum),
    .io_in_flow(PE_Array_21_8_io_in_flow),
    .io_in_shift(PE_Array_21_8_io_in_shift),
    .io_out_activate(PE_Array_21_8_io_out_activate),
    .io_out_weight(PE_Array_21_8_io_out_weight),
    .io_out_psum(PE_Array_21_8_io_out_psum)
  );
  basic_PE PE_Array_21_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_9_clock),
    .reset(PE_Array_21_9_reset),
    .io_in_activate(PE_Array_21_9_io_in_activate),
    .io_in_weight(PE_Array_21_9_io_in_weight),
    .io_in_psum(PE_Array_21_9_io_in_psum),
    .io_in_flow(PE_Array_21_9_io_in_flow),
    .io_in_shift(PE_Array_21_9_io_in_shift),
    .io_out_activate(PE_Array_21_9_io_out_activate),
    .io_out_weight(PE_Array_21_9_io_out_weight),
    .io_out_psum(PE_Array_21_9_io_out_psum)
  );
  basic_PE PE_Array_21_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_10_clock),
    .reset(PE_Array_21_10_reset),
    .io_in_activate(PE_Array_21_10_io_in_activate),
    .io_in_weight(PE_Array_21_10_io_in_weight),
    .io_in_psum(PE_Array_21_10_io_in_psum),
    .io_in_flow(PE_Array_21_10_io_in_flow),
    .io_in_shift(PE_Array_21_10_io_in_shift),
    .io_out_activate(PE_Array_21_10_io_out_activate),
    .io_out_weight(PE_Array_21_10_io_out_weight),
    .io_out_psum(PE_Array_21_10_io_out_psum)
  );
  basic_PE PE_Array_21_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_11_clock),
    .reset(PE_Array_21_11_reset),
    .io_in_activate(PE_Array_21_11_io_in_activate),
    .io_in_weight(PE_Array_21_11_io_in_weight),
    .io_in_psum(PE_Array_21_11_io_in_psum),
    .io_in_flow(PE_Array_21_11_io_in_flow),
    .io_in_shift(PE_Array_21_11_io_in_shift),
    .io_out_activate(PE_Array_21_11_io_out_activate),
    .io_out_weight(PE_Array_21_11_io_out_weight),
    .io_out_psum(PE_Array_21_11_io_out_psum)
  );
  basic_PE PE_Array_21_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_12_clock),
    .reset(PE_Array_21_12_reset),
    .io_in_activate(PE_Array_21_12_io_in_activate),
    .io_in_weight(PE_Array_21_12_io_in_weight),
    .io_in_psum(PE_Array_21_12_io_in_psum),
    .io_in_flow(PE_Array_21_12_io_in_flow),
    .io_in_shift(PE_Array_21_12_io_in_shift),
    .io_out_activate(PE_Array_21_12_io_out_activate),
    .io_out_weight(PE_Array_21_12_io_out_weight),
    .io_out_psum(PE_Array_21_12_io_out_psum)
  );
  basic_PE PE_Array_21_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_13_clock),
    .reset(PE_Array_21_13_reset),
    .io_in_activate(PE_Array_21_13_io_in_activate),
    .io_in_weight(PE_Array_21_13_io_in_weight),
    .io_in_psum(PE_Array_21_13_io_in_psum),
    .io_in_flow(PE_Array_21_13_io_in_flow),
    .io_in_shift(PE_Array_21_13_io_in_shift),
    .io_out_activate(PE_Array_21_13_io_out_activate),
    .io_out_weight(PE_Array_21_13_io_out_weight),
    .io_out_psum(PE_Array_21_13_io_out_psum)
  );
  basic_PE PE_Array_21_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_14_clock),
    .reset(PE_Array_21_14_reset),
    .io_in_activate(PE_Array_21_14_io_in_activate),
    .io_in_weight(PE_Array_21_14_io_in_weight),
    .io_in_psum(PE_Array_21_14_io_in_psum),
    .io_in_flow(PE_Array_21_14_io_in_flow),
    .io_in_shift(PE_Array_21_14_io_in_shift),
    .io_out_activate(PE_Array_21_14_io_out_activate),
    .io_out_weight(PE_Array_21_14_io_out_weight),
    .io_out_psum(PE_Array_21_14_io_out_psum)
  );
  basic_PE PE_Array_21_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_15_clock),
    .reset(PE_Array_21_15_reset),
    .io_in_activate(PE_Array_21_15_io_in_activate),
    .io_in_weight(PE_Array_21_15_io_in_weight),
    .io_in_psum(PE_Array_21_15_io_in_psum),
    .io_in_flow(PE_Array_21_15_io_in_flow),
    .io_in_shift(PE_Array_21_15_io_in_shift),
    .io_out_activate(PE_Array_21_15_io_out_activate),
    .io_out_weight(PE_Array_21_15_io_out_weight),
    .io_out_psum(PE_Array_21_15_io_out_psum)
  );
  basic_PE PE_Array_21_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_16_clock),
    .reset(PE_Array_21_16_reset),
    .io_in_activate(PE_Array_21_16_io_in_activate),
    .io_in_weight(PE_Array_21_16_io_in_weight),
    .io_in_psum(PE_Array_21_16_io_in_psum),
    .io_in_flow(PE_Array_21_16_io_in_flow),
    .io_in_shift(PE_Array_21_16_io_in_shift),
    .io_out_activate(PE_Array_21_16_io_out_activate),
    .io_out_weight(PE_Array_21_16_io_out_weight),
    .io_out_psum(PE_Array_21_16_io_out_psum)
  );
  basic_PE PE_Array_21_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_17_clock),
    .reset(PE_Array_21_17_reset),
    .io_in_activate(PE_Array_21_17_io_in_activate),
    .io_in_weight(PE_Array_21_17_io_in_weight),
    .io_in_psum(PE_Array_21_17_io_in_psum),
    .io_in_flow(PE_Array_21_17_io_in_flow),
    .io_in_shift(PE_Array_21_17_io_in_shift),
    .io_out_activate(PE_Array_21_17_io_out_activate),
    .io_out_weight(PE_Array_21_17_io_out_weight),
    .io_out_psum(PE_Array_21_17_io_out_psum)
  );
  basic_PE PE_Array_21_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_18_clock),
    .reset(PE_Array_21_18_reset),
    .io_in_activate(PE_Array_21_18_io_in_activate),
    .io_in_weight(PE_Array_21_18_io_in_weight),
    .io_in_psum(PE_Array_21_18_io_in_psum),
    .io_in_flow(PE_Array_21_18_io_in_flow),
    .io_in_shift(PE_Array_21_18_io_in_shift),
    .io_out_activate(PE_Array_21_18_io_out_activate),
    .io_out_weight(PE_Array_21_18_io_out_weight),
    .io_out_psum(PE_Array_21_18_io_out_psum)
  );
  basic_PE PE_Array_21_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_19_clock),
    .reset(PE_Array_21_19_reset),
    .io_in_activate(PE_Array_21_19_io_in_activate),
    .io_in_weight(PE_Array_21_19_io_in_weight),
    .io_in_psum(PE_Array_21_19_io_in_psum),
    .io_in_flow(PE_Array_21_19_io_in_flow),
    .io_in_shift(PE_Array_21_19_io_in_shift),
    .io_out_activate(PE_Array_21_19_io_out_activate),
    .io_out_weight(PE_Array_21_19_io_out_weight),
    .io_out_psum(PE_Array_21_19_io_out_psum)
  );
  basic_PE PE_Array_21_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_20_clock),
    .reset(PE_Array_21_20_reset),
    .io_in_activate(PE_Array_21_20_io_in_activate),
    .io_in_weight(PE_Array_21_20_io_in_weight),
    .io_in_psum(PE_Array_21_20_io_in_psum),
    .io_in_flow(PE_Array_21_20_io_in_flow),
    .io_in_shift(PE_Array_21_20_io_in_shift),
    .io_out_activate(PE_Array_21_20_io_out_activate),
    .io_out_weight(PE_Array_21_20_io_out_weight),
    .io_out_psum(PE_Array_21_20_io_out_psum)
  );
  basic_PE PE_Array_21_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_21_clock),
    .reset(PE_Array_21_21_reset),
    .io_in_activate(PE_Array_21_21_io_in_activate),
    .io_in_weight(PE_Array_21_21_io_in_weight),
    .io_in_psum(PE_Array_21_21_io_in_psum),
    .io_in_flow(PE_Array_21_21_io_in_flow),
    .io_in_shift(PE_Array_21_21_io_in_shift),
    .io_out_activate(PE_Array_21_21_io_out_activate),
    .io_out_weight(PE_Array_21_21_io_out_weight),
    .io_out_psum(PE_Array_21_21_io_out_psum)
  );
  basic_PE PE_Array_21_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_22_clock),
    .reset(PE_Array_21_22_reset),
    .io_in_activate(PE_Array_21_22_io_in_activate),
    .io_in_weight(PE_Array_21_22_io_in_weight),
    .io_in_psum(PE_Array_21_22_io_in_psum),
    .io_in_flow(PE_Array_21_22_io_in_flow),
    .io_in_shift(PE_Array_21_22_io_in_shift),
    .io_out_activate(PE_Array_21_22_io_out_activate),
    .io_out_weight(PE_Array_21_22_io_out_weight),
    .io_out_psum(PE_Array_21_22_io_out_psum)
  );
  basic_PE PE_Array_21_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_23_clock),
    .reset(PE_Array_21_23_reset),
    .io_in_activate(PE_Array_21_23_io_in_activate),
    .io_in_weight(PE_Array_21_23_io_in_weight),
    .io_in_psum(PE_Array_21_23_io_in_psum),
    .io_in_flow(PE_Array_21_23_io_in_flow),
    .io_in_shift(PE_Array_21_23_io_in_shift),
    .io_out_activate(PE_Array_21_23_io_out_activate),
    .io_out_weight(PE_Array_21_23_io_out_weight),
    .io_out_psum(PE_Array_21_23_io_out_psum)
  );
  basic_PE PE_Array_21_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_24_clock),
    .reset(PE_Array_21_24_reset),
    .io_in_activate(PE_Array_21_24_io_in_activate),
    .io_in_weight(PE_Array_21_24_io_in_weight),
    .io_in_psum(PE_Array_21_24_io_in_psum),
    .io_in_flow(PE_Array_21_24_io_in_flow),
    .io_in_shift(PE_Array_21_24_io_in_shift),
    .io_out_activate(PE_Array_21_24_io_out_activate),
    .io_out_weight(PE_Array_21_24_io_out_weight),
    .io_out_psum(PE_Array_21_24_io_out_psum)
  );
  basic_PE PE_Array_21_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_25_clock),
    .reset(PE_Array_21_25_reset),
    .io_in_activate(PE_Array_21_25_io_in_activate),
    .io_in_weight(PE_Array_21_25_io_in_weight),
    .io_in_psum(PE_Array_21_25_io_in_psum),
    .io_in_flow(PE_Array_21_25_io_in_flow),
    .io_in_shift(PE_Array_21_25_io_in_shift),
    .io_out_activate(PE_Array_21_25_io_out_activate),
    .io_out_weight(PE_Array_21_25_io_out_weight),
    .io_out_psum(PE_Array_21_25_io_out_psum)
  );
  basic_PE PE_Array_21_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_26_clock),
    .reset(PE_Array_21_26_reset),
    .io_in_activate(PE_Array_21_26_io_in_activate),
    .io_in_weight(PE_Array_21_26_io_in_weight),
    .io_in_psum(PE_Array_21_26_io_in_psum),
    .io_in_flow(PE_Array_21_26_io_in_flow),
    .io_in_shift(PE_Array_21_26_io_in_shift),
    .io_out_activate(PE_Array_21_26_io_out_activate),
    .io_out_weight(PE_Array_21_26_io_out_weight),
    .io_out_psum(PE_Array_21_26_io_out_psum)
  );
  basic_PE PE_Array_21_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_27_clock),
    .reset(PE_Array_21_27_reset),
    .io_in_activate(PE_Array_21_27_io_in_activate),
    .io_in_weight(PE_Array_21_27_io_in_weight),
    .io_in_psum(PE_Array_21_27_io_in_psum),
    .io_in_flow(PE_Array_21_27_io_in_flow),
    .io_in_shift(PE_Array_21_27_io_in_shift),
    .io_out_activate(PE_Array_21_27_io_out_activate),
    .io_out_weight(PE_Array_21_27_io_out_weight),
    .io_out_psum(PE_Array_21_27_io_out_psum)
  );
  basic_PE PE_Array_21_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_28_clock),
    .reset(PE_Array_21_28_reset),
    .io_in_activate(PE_Array_21_28_io_in_activate),
    .io_in_weight(PE_Array_21_28_io_in_weight),
    .io_in_psum(PE_Array_21_28_io_in_psum),
    .io_in_flow(PE_Array_21_28_io_in_flow),
    .io_in_shift(PE_Array_21_28_io_in_shift),
    .io_out_activate(PE_Array_21_28_io_out_activate),
    .io_out_weight(PE_Array_21_28_io_out_weight),
    .io_out_psum(PE_Array_21_28_io_out_psum)
  );
  basic_PE PE_Array_21_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_29_clock),
    .reset(PE_Array_21_29_reset),
    .io_in_activate(PE_Array_21_29_io_in_activate),
    .io_in_weight(PE_Array_21_29_io_in_weight),
    .io_in_psum(PE_Array_21_29_io_in_psum),
    .io_in_flow(PE_Array_21_29_io_in_flow),
    .io_in_shift(PE_Array_21_29_io_in_shift),
    .io_out_activate(PE_Array_21_29_io_out_activate),
    .io_out_weight(PE_Array_21_29_io_out_weight),
    .io_out_psum(PE_Array_21_29_io_out_psum)
  );
  basic_PE PE_Array_21_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_30_clock),
    .reset(PE_Array_21_30_reset),
    .io_in_activate(PE_Array_21_30_io_in_activate),
    .io_in_weight(PE_Array_21_30_io_in_weight),
    .io_in_psum(PE_Array_21_30_io_in_psum),
    .io_in_flow(PE_Array_21_30_io_in_flow),
    .io_in_shift(PE_Array_21_30_io_in_shift),
    .io_out_activate(PE_Array_21_30_io_out_activate),
    .io_out_weight(PE_Array_21_30_io_out_weight),
    .io_out_psum(PE_Array_21_30_io_out_psum)
  );
  basic_PE PE_Array_21_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_21_31_clock),
    .reset(PE_Array_21_31_reset),
    .io_in_activate(PE_Array_21_31_io_in_activate),
    .io_in_weight(PE_Array_21_31_io_in_weight),
    .io_in_psum(PE_Array_21_31_io_in_psum),
    .io_in_flow(PE_Array_21_31_io_in_flow),
    .io_in_shift(PE_Array_21_31_io_in_shift),
    .io_out_activate(PE_Array_21_31_io_out_activate),
    .io_out_weight(PE_Array_21_31_io_out_weight),
    .io_out_psum(PE_Array_21_31_io_out_psum)
  );
  basic_PE PE_Array_22_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_0_clock),
    .reset(PE_Array_22_0_reset),
    .io_in_activate(PE_Array_22_0_io_in_activate),
    .io_in_weight(PE_Array_22_0_io_in_weight),
    .io_in_psum(PE_Array_22_0_io_in_psum),
    .io_in_flow(PE_Array_22_0_io_in_flow),
    .io_in_shift(PE_Array_22_0_io_in_shift),
    .io_out_activate(PE_Array_22_0_io_out_activate),
    .io_out_weight(PE_Array_22_0_io_out_weight),
    .io_out_psum(PE_Array_22_0_io_out_psum)
  );
  basic_PE PE_Array_22_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_1_clock),
    .reset(PE_Array_22_1_reset),
    .io_in_activate(PE_Array_22_1_io_in_activate),
    .io_in_weight(PE_Array_22_1_io_in_weight),
    .io_in_psum(PE_Array_22_1_io_in_psum),
    .io_in_flow(PE_Array_22_1_io_in_flow),
    .io_in_shift(PE_Array_22_1_io_in_shift),
    .io_out_activate(PE_Array_22_1_io_out_activate),
    .io_out_weight(PE_Array_22_1_io_out_weight),
    .io_out_psum(PE_Array_22_1_io_out_psum)
  );
  basic_PE PE_Array_22_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_2_clock),
    .reset(PE_Array_22_2_reset),
    .io_in_activate(PE_Array_22_2_io_in_activate),
    .io_in_weight(PE_Array_22_2_io_in_weight),
    .io_in_psum(PE_Array_22_2_io_in_psum),
    .io_in_flow(PE_Array_22_2_io_in_flow),
    .io_in_shift(PE_Array_22_2_io_in_shift),
    .io_out_activate(PE_Array_22_2_io_out_activate),
    .io_out_weight(PE_Array_22_2_io_out_weight),
    .io_out_psum(PE_Array_22_2_io_out_psum)
  );
  basic_PE PE_Array_22_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_3_clock),
    .reset(PE_Array_22_3_reset),
    .io_in_activate(PE_Array_22_3_io_in_activate),
    .io_in_weight(PE_Array_22_3_io_in_weight),
    .io_in_psum(PE_Array_22_3_io_in_psum),
    .io_in_flow(PE_Array_22_3_io_in_flow),
    .io_in_shift(PE_Array_22_3_io_in_shift),
    .io_out_activate(PE_Array_22_3_io_out_activate),
    .io_out_weight(PE_Array_22_3_io_out_weight),
    .io_out_psum(PE_Array_22_3_io_out_psum)
  );
  basic_PE PE_Array_22_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_4_clock),
    .reset(PE_Array_22_4_reset),
    .io_in_activate(PE_Array_22_4_io_in_activate),
    .io_in_weight(PE_Array_22_4_io_in_weight),
    .io_in_psum(PE_Array_22_4_io_in_psum),
    .io_in_flow(PE_Array_22_4_io_in_flow),
    .io_in_shift(PE_Array_22_4_io_in_shift),
    .io_out_activate(PE_Array_22_4_io_out_activate),
    .io_out_weight(PE_Array_22_4_io_out_weight),
    .io_out_psum(PE_Array_22_4_io_out_psum)
  );
  basic_PE PE_Array_22_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_5_clock),
    .reset(PE_Array_22_5_reset),
    .io_in_activate(PE_Array_22_5_io_in_activate),
    .io_in_weight(PE_Array_22_5_io_in_weight),
    .io_in_psum(PE_Array_22_5_io_in_psum),
    .io_in_flow(PE_Array_22_5_io_in_flow),
    .io_in_shift(PE_Array_22_5_io_in_shift),
    .io_out_activate(PE_Array_22_5_io_out_activate),
    .io_out_weight(PE_Array_22_5_io_out_weight),
    .io_out_psum(PE_Array_22_5_io_out_psum)
  );
  basic_PE PE_Array_22_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_6_clock),
    .reset(PE_Array_22_6_reset),
    .io_in_activate(PE_Array_22_6_io_in_activate),
    .io_in_weight(PE_Array_22_6_io_in_weight),
    .io_in_psum(PE_Array_22_6_io_in_psum),
    .io_in_flow(PE_Array_22_6_io_in_flow),
    .io_in_shift(PE_Array_22_6_io_in_shift),
    .io_out_activate(PE_Array_22_6_io_out_activate),
    .io_out_weight(PE_Array_22_6_io_out_weight),
    .io_out_psum(PE_Array_22_6_io_out_psum)
  );
  basic_PE PE_Array_22_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_7_clock),
    .reset(PE_Array_22_7_reset),
    .io_in_activate(PE_Array_22_7_io_in_activate),
    .io_in_weight(PE_Array_22_7_io_in_weight),
    .io_in_psum(PE_Array_22_7_io_in_psum),
    .io_in_flow(PE_Array_22_7_io_in_flow),
    .io_in_shift(PE_Array_22_7_io_in_shift),
    .io_out_activate(PE_Array_22_7_io_out_activate),
    .io_out_weight(PE_Array_22_7_io_out_weight),
    .io_out_psum(PE_Array_22_7_io_out_psum)
  );
  basic_PE PE_Array_22_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_8_clock),
    .reset(PE_Array_22_8_reset),
    .io_in_activate(PE_Array_22_8_io_in_activate),
    .io_in_weight(PE_Array_22_8_io_in_weight),
    .io_in_psum(PE_Array_22_8_io_in_psum),
    .io_in_flow(PE_Array_22_8_io_in_flow),
    .io_in_shift(PE_Array_22_8_io_in_shift),
    .io_out_activate(PE_Array_22_8_io_out_activate),
    .io_out_weight(PE_Array_22_8_io_out_weight),
    .io_out_psum(PE_Array_22_8_io_out_psum)
  );
  basic_PE PE_Array_22_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_9_clock),
    .reset(PE_Array_22_9_reset),
    .io_in_activate(PE_Array_22_9_io_in_activate),
    .io_in_weight(PE_Array_22_9_io_in_weight),
    .io_in_psum(PE_Array_22_9_io_in_psum),
    .io_in_flow(PE_Array_22_9_io_in_flow),
    .io_in_shift(PE_Array_22_9_io_in_shift),
    .io_out_activate(PE_Array_22_9_io_out_activate),
    .io_out_weight(PE_Array_22_9_io_out_weight),
    .io_out_psum(PE_Array_22_9_io_out_psum)
  );
  basic_PE PE_Array_22_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_10_clock),
    .reset(PE_Array_22_10_reset),
    .io_in_activate(PE_Array_22_10_io_in_activate),
    .io_in_weight(PE_Array_22_10_io_in_weight),
    .io_in_psum(PE_Array_22_10_io_in_psum),
    .io_in_flow(PE_Array_22_10_io_in_flow),
    .io_in_shift(PE_Array_22_10_io_in_shift),
    .io_out_activate(PE_Array_22_10_io_out_activate),
    .io_out_weight(PE_Array_22_10_io_out_weight),
    .io_out_psum(PE_Array_22_10_io_out_psum)
  );
  basic_PE PE_Array_22_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_11_clock),
    .reset(PE_Array_22_11_reset),
    .io_in_activate(PE_Array_22_11_io_in_activate),
    .io_in_weight(PE_Array_22_11_io_in_weight),
    .io_in_psum(PE_Array_22_11_io_in_psum),
    .io_in_flow(PE_Array_22_11_io_in_flow),
    .io_in_shift(PE_Array_22_11_io_in_shift),
    .io_out_activate(PE_Array_22_11_io_out_activate),
    .io_out_weight(PE_Array_22_11_io_out_weight),
    .io_out_psum(PE_Array_22_11_io_out_psum)
  );
  basic_PE PE_Array_22_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_12_clock),
    .reset(PE_Array_22_12_reset),
    .io_in_activate(PE_Array_22_12_io_in_activate),
    .io_in_weight(PE_Array_22_12_io_in_weight),
    .io_in_psum(PE_Array_22_12_io_in_psum),
    .io_in_flow(PE_Array_22_12_io_in_flow),
    .io_in_shift(PE_Array_22_12_io_in_shift),
    .io_out_activate(PE_Array_22_12_io_out_activate),
    .io_out_weight(PE_Array_22_12_io_out_weight),
    .io_out_psum(PE_Array_22_12_io_out_psum)
  );
  basic_PE PE_Array_22_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_13_clock),
    .reset(PE_Array_22_13_reset),
    .io_in_activate(PE_Array_22_13_io_in_activate),
    .io_in_weight(PE_Array_22_13_io_in_weight),
    .io_in_psum(PE_Array_22_13_io_in_psum),
    .io_in_flow(PE_Array_22_13_io_in_flow),
    .io_in_shift(PE_Array_22_13_io_in_shift),
    .io_out_activate(PE_Array_22_13_io_out_activate),
    .io_out_weight(PE_Array_22_13_io_out_weight),
    .io_out_psum(PE_Array_22_13_io_out_psum)
  );
  basic_PE PE_Array_22_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_14_clock),
    .reset(PE_Array_22_14_reset),
    .io_in_activate(PE_Array_22_14_io_in_activate),
    .io_in_weight(PE_Array_22_14_io_in_weight),
    .io_in_psum(PE_Array_22_14_io_in_psum),
    .io_in_flow(PE_Array_22_14_io_in_flow),
    .io_in_shift(PE_Array_22_14_io_in_shift),
    .io_out_activate(PE_Array_22_14_io_out_activate),
    .io_out_weight(PE_Array_22_14_io_out_weight),
    .io_out_psum(PE_Array_22_14_io_out_psum)
  );
  basic_PE PE_Array_22_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_15_clock),
    .reset(PE_Array_22_15_reset),
    .io_in_activate(PE_Array_22_15_io_in_activate),
    .io_in_weight(PE_Array_22_15_io_in_weight),
    .io_in_psum(PE_Array_22_15_io_in_psum),
    .io_in_flow(PE_Array_22_15_io_in_flow),
    .io_in_shift(PE_Array_22_15_io_in_shift),
    .io_out_activate(PE_Array_22_15_io_out_activate),
    .io_out_weight(PE_Array_22_15_io_out_weight),
    .io_out_psum(PE_Array_22_15_io_out_psum)
  );
  basic_PE PE_Array_22_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_16_clock),
    .reset(PE_Array_22_16_reset),
    .io_in_activate(PE_Array_22_16_io_in_activate),
    .io_in_weight(PE_Array_22_16_io_in_weight),
    .io_in_psum(PE_Array_22_16_io_in_psum),
    .io_in_flow(PE_Array_22_16_io_in_flow),
    .io_in_shift(PE_Array_22_16_io_in_shift),
    .io_out_activate(PE_Array_22_16_io_out_activate),
    .io_out_weight(PE_Array_22_16_io_out_weight),
    .io_out_psum(PE_Array_22_16_io_out_psum)
  );
  basic_PE PE_Array_22_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_17_clock),
    .reset(PE_Array_22_17_reset),
    .io_in_activate(PE_Array_22_17_io_in_activate),
    .io_in_weight(PE_Array_22_17_io_in_weight),
    .io_in_psum(PE_Array_22_17_io_in_psum),
    .io_in_flow(PE_Array_22_17_io_in_flow),
    .io_in_shift(PE_Array_22_17_io_in_shift),
    .io_out_activate(PE_Array_22_17_io_out_activate),
    .io_out_weight(PE_Array_22_17_io_out_weight),
    .io_out_psum(PE_Array_22_17_io_out_psum)
  );
  basic_PE PE_Array_22_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_18_clock),
    .reset(PE_Array_22_18_reset),
    .io_in_activate(PE_Array_22_18_io_in_activate),
    .io_in_weight(PE_Array_22_18_io_in_weight),
    .io_in_psum(PE_Array_22_18_io_in_psum),
    .io_in_flow(PE_Array_22_18_io_in_flow),
    .io_in_shift(PE_Array_22_18_io_in_shift),
    .io_out_activate(PE_Array_22_18_io_out_activate),
    .io_out_weight(PE_Array_22_18_io_out_weight),
    .io_out_psum(PE_Array_22_18_io_out_psum)
  );
  basic_PE PE_Array_22_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_19_clock),
    .reset(PE_Array_22_19_reset),
    .io_in_activate(PE_Array_22_19_io_in_activate),
    .io_in_weight(PE_Array_22_19_io_in_weight),
    .io_in_psum(PE_Array_22_19_io_in_psum),
    .io_in_flow(PE_Array_22_19_io_in_flow),
    .io_in_shift(PE_Array_22_19_io_in_shift),
    .io_out_activate(PE_Array_22_19_io_out_activate),
    .io_out_weight(PE_Array_22_19_io_out_weight),
    .io_out_psum(PE_Array_22_19_io_out_psum)
  );
  basic_PE PE_Array_22_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_20_clock),
    .reset(PE_Array_22_20_reset),
    .io_in_activate(PE_Array_22_20_io_in_activate),
    .io_in_weight(PE_Array_22_20_io_in_weight),
    .io_in_psum(PE_Array_22_20_io_in_psum),
    .io_in_flow(PE_Array_22_20_io_in_flow),
    .io_in_shift(PE_Array_22_20_io_in_shift),
    .io_out_activate(PE_Array_22_20_io_out_activate),
    .io_out_weight(PE_Array_22_20_io_out_weight),
    .io_out_psum(PE_Array_22_20_io_out_psum)
  );
  basic_PE PE_Array_22_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_21_clock),
    .reset(PE_Array_22_21_reset),
    .io_in_activate(PE_Array_22_21_io_in_activate),
    .io_in_weight(PE_Array_22_21_io_in_weight),
    .io_in_psum(PE_Array_22_21_io_in_psum),
    .io_in_flow(PE_Array_22_21_io_in_flow),
    .io_in_shift(PE_Array_22_21_io_in_shift),
    .io_out_activate(PE_Array_22_21_io_out_activate),
    .io_out_weight(PE_Array_22_21_io_out_weight),
    .io_out_psum(PE_Array_22_21_io_out_psum)
  );
  basic_PE PE_Array_22_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_22_clock),
    .reset(PE_Array_22_22_reset),
    .io_in_activate(PE_Array_22_22_io_in_activate),
    .io_in_weight(PE_Array_22_22_io_in_weight),
    .io_in_psum(PE_Array_22_22_io_in_psum),
    .io_in_flow(PE_Array_22_22_io_in_flow),
    .io_in_shift(PE_Array_22_22_io_in_shift),
    .io_out_activate(PE_Array_22_22_io_out_activate),
    .io_out_weight(PE_Array_22_22_io_out_weight),
    .io_out_psum(PE_Array_22_22_io_out_psum)
  );
  basic_PE PE_Array_22_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_23_clock),
    .reset(PE_Array_22_23_reset),
    .io_in_activate(PE_Array_22_23_io_in_activate),
    .io_in_weight(PE_Array_22_23_io_in_weight),
    .io_in_psum(PE_Array_22_23_io_in_psum),
    .io_in_flow(PE_Array_22_23_io_in_flow),
    .io_in_shift(PE_Array_22_23_io_in_shift),
    .io_out_activate(PE_Array_22_23_io_out_activate),
    .io_out_weight(PE_Array_22_23_io_out_weight),
    .io_out_psum(PE_Array_22_23_io_out_psum)
  );
  basic_PE PE_Array_22_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_24_clock),
    .reset(PE_Array_22_24_reset),
    .io_in_activate(PE_Array_22_24_io_in_activate),
    .io_in_weight(PE_Array_22_24_io_in_weight),
    .io_in_psum(PE_Array_22_24_io_in_psum),
    .io_in_flow(PE_Array_22_24_io_in_flow),
    .io_in_shift(PE_Array_22_24_io_in_shift),
    .io_out_activate(PE_Array_22_24_io_out_activate),
    .io_out_weight(PE_Array_22_24_io_out_weight),
    .io_out_psum(PE_Array_22_24_io_out_psum)
  );
  basic_PE PE_Array_22_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_25_clock),
    .reset(PE_Array_22_25_reset),
    .io_in_activate(PE_Array_22_25_io_in_activate),
    .io_in_weight(PE_Array_22_25_io_in_weight),
    .io_in_psum(PE_Array_22_25_io_in_psum),
    .io_in_flow(PE_Array_22_25_io_in_flow),
    .io_in_shift(PE_Array_22_25_io_in_shift),
    .io_out_activate(PE_Array_22_25_io_out_activate),
    .io_out_weight(PE_Array_22_25_io_out_weight),
    .io_out_psum(PE_Array_22_25_io_out_psum)
  );
  basic_PE PE_Array_22_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_26_clock),
    .reset(PE_Array_22_26_reset),
    .io_in_activate(PE_Array_22_26_io_in_activate),
    .io_in_weight(PE_Array_22_26_io_in_weight),
    .io_in_psum(PE_Array_22_26_io_in_psum),
    .io_in_flow(PE_Array_22_26_io_in_flow),
    .io_in_shift(PE_Array_22_26_io_in_shift),
    .io_out_activate(PE_Array_22_26_io_out_activate),
    .io_out_weight(PE_Array_22_26_io_out_weight),
    .io_out_psum(PE_Array_22_26_io_out_psum)
  );
  basic_PE PE_Array_22_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_27_clock),
    .reset(PE_Array_22_27_reset),
    .io_in_activate(PE_Array_22_27_io_in_activate),
    .io_in_weight(PE_Array_22_27_io_in_weight),
    .io_in_psum(PE_Array_22_27_io_in_psum),
    .io_in_flow(PE_Array_22_27_io_in_flow),
    .io_in_shift(PE_Array_22_27_io_in_shift),
    .io_out_activate(PE_Array_22_27_io_out_activate),
    .io_out_weight(PE_Array_22_27_io_out_weight),
    .io_out_psum(PE_Array_22_27_io_out_psum)
  );
  basic_PE PE_Array_22_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_28_clock),
    .reset(PE_Array_22_28_reset),
    .io_in_activate(PE_Array_22_28_io_in_activate),
    .io_in_weight(PE_Array_22_28_io_in_weight),
    .io_in_psum(PE_Array_22_28_io_in_psum),
    .io_in_flow(PE_Array_22_28_io_in_flow),
    .io_in_shift(PE_Array_22_28_io_in_shift),
    .io_out_activate(PE_Array_22_28_io_out_activate),
    .io_out_weight(PE_Array_22_28_io_out_weight),
    .io_out_psum(PE_Array_22_28_io_out_psum)
  );
  basic_PE PE_Array_22_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_29_clock),
    .reset(PE_Array_22_29_reset),
    .io_in_activate(PE_Array_22_29_io_in_activate),
    .io_in_weight(PE_Array_22_29_io_in_weight),
    .io_in_psum(PE_Array_22_29_io_in_psum),
    .io_in_flow(PE_Array_22_29_io_in_flow),
    .io_in_shift(PE_Array_22_29_io_in_shift),
    .io_out_activate(PE_Array_22_29_io_out_activate),
    .io_out_weight(PE_Array_22_29_io_out_weight),
    .io_out_psum(PE_Array_22_29_io_out_psum)
  );
  basic_PE PE_Array_22_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_30_clock),
    .reset(PE_Array_22_30_reset),
    .io_in_activate(PE_Array_22_30_io_in_activate),
    .io_in_weight(PE_Array_22_30_io_in_weight),
    .io_in_psum(PE_Array_22_30_io_in_psum),
    .io_in_flow(PE_Array_22_30_io_in_flow),
    .io_in_shift(PE_Array_22_30_io_in_shift),
    .io_out_activate(PE_Array_22_30_io_out_activate),
    .io_out_weight(PE_Array_22_30_io_out_weight),
    .io_out_psum(PE_Array_22_30_io_out_psum)
  );
  basic_PE PE_Array_22_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_22_31_clock),
    .reset(PE_Array_22_31_reset),
    .io_in_activate(PE_Array_22_31_io_in_activate),
    .io_in_weight(PE_Array_22_31_io_in_weight),
    .io_in_psum(PE_Array_22_31_io_in_psum),
    .io_in_flow(PE_Array_22_31_io_in_flow),
    .io_in_shift(PE_Array_22_31_io_in_shift),
    .io_out_activate(PE_Array_22_31_io_out_activate),
    .io_out_weight(PE_Array_22_31_io_out_weight),
    .io_out_psum(PE_Array_22_31_io_out_psum)
  );
  basic_PE PE_Array_23_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_0_clock),
    .reset(PE_Array_23_0_reset),
    .io_in_activate(PE_Array_23_0_io_in_activate),
    .io_in_weight(PE_Array_23_0_io_in_weight),
    .io_in_psum(PE_Array_23_0_io_in_psum),
    .io_in_flow(PE_Array_23_0_io_in_flow),
    .io_in_shift(PE_Array_23_0_io_in_shift),
    .io_out_activate(PE_Array_23_0_io_out_activate),
    .io_out_weight(PE_Array_23_0_io_out_weight),
    .io_out_psum(PE_Array_23_0_io_out_psum)
  );
  basic_PE PE_Array_23_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_1_clock),
    .reset(PE_Array_23_1_reset),
    .io_in_activate(PE_Array_23_1_io_in_activate),
    .io_in_weight(PE_Array_23_1_io_in_weight),
    .io_in_psum(PE_Array_23_1_io_in_psum),
    .io_in_flow(PE_Array_23_1_io_in_flow),
    .io_in_shift(PE_Array_23_1_io_in_shift),
    .io_out_activate(PE_Array_23_1_io_out_activate),
    .io_out_weight(PE_Array_23_1_io_out_weight),
    .io_out_psum(PE_Array_23_1_io_out_psum)
  );
  basic_PE PE_Array_23_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_2_clock),
    .reset(PE_Array_23_2_reset),
    .io_in_activate(PE_Array_23_2_io_in_activate),
    .io_in_weight(PE_Array_23_2_io_in_weight),
    .io_in_psum(PE_Array_23_2_io_in_psum),
    .io_in_flow(PE_Array_23_2_io_in_flow),
    .io_in_shift(PE_Array_23_2_io_in_shift),
    .io_out_activate(PE_Array_23_2_io_out_activate),
    .io_out_weight(PE_Array_23_2_io_out_weight),
    .io_out_psum(PE_Array_23_2_io_out_psum)
  );
  basic_PE PE_Array_23_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_3_clock),
    .reset(PE_Array_23_3_reset),
    .io_in_activate(PE_Array_23_3_io_in_activate),
    .io_in_weight(PE_Array_23_3_io_in_weight),
    .io_in_psum(PE_Array_23_3_io_in_psum),
    .io_in_flow(PE_Array_23_3_io_in_flow),
    .io_in_shift(PE_Array_23_3_io_in_shift),
    .io_out_activate(PE_Array_23_3_io_out_activate),
    .io_out_weight(PE_Array_23_3_io_out_weight),
    .io_out_psum(PE_Array_23_3_io_out_psum)
  );
  basic_PE PE_Array_23_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_4_clock),
    .reset(PE_Array_23_4_reset),
    .io_in_activate(PE_Array_23_4_io_in_activate),
    .io_in_weight(PE_Array_23_4_io_in_weight),
    .io_in_psum(PE_Array_23_4_io_in_psum),
    .io_in_flow(PE_Array_23_4_io_in_flow),
    .io_in_shift(PE_Array_23_4_io_in_shift),
    .io_out_activate(PE_Array_23_4_io_out_activate),
    .io_out_weight(PE_Array_23_4_io_out_weight),
    .io_out_psum(PE_Array_23_4_io_out_psum)
  );
  basic_PE PE_Array_23_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_5_clock),
    .reset(PE_Array_23_5_reset),
    .io_in_activate(PE_Array_23_5_io_in_activate),
    .io_in_weight(PE_Array_23_5_io_in_weight),
    .io_in_psum(PE_Array_23_5_io_in_psum),
    .io_in_flow(PE_Array_23_5_io_in_flow),
    .io_in_shift(PE_Array_23_5_io_in_shift),
    .io_out_activate(PE_Array_23_5_io_out_activate),
    .io_out_weight(PE_Array_23_5_io_out_weight),
    .io_out_psum(PE_Array_23_5_io_out_psum)
  );
  basic_PE PE_Array_23_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_6_clock),
    .reset(PE_Array_23_6_reset),
    .io_in_activate(PE_Array_23_6_io_in_activate),
    .io_in_weight(PE_Array_23_6_io_in_weight),
    .io_in_psum(PE_Array_23_6_io_in_psum),
    .io_in_flow(PE_Array_23_6_io_in_flow),
    .io_in_shift(PE_Array_23_6_io_in_shift),
    .io_out_activate(PE_Array_23_6_io_out_activate),
    .io_out_weight(PE_Array_23_6_io_out_weight),
    .io_out_psum(PE_Array_23_6_io_out_psum)
  );
  basic_PE PE_Array_23_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_7_clock),
    .reset(PE_Array_23_7_reset),
    .io_in_activate(PE_Array_23_7_io_in_activate),
    .io_in_weight(PE_Array_23_7_io_in_weight),
    .io_in_psum(PE_Array_23_7_io_in_psum),
    .io_in_flow(PE_Array_23_7_io_in_flow),
    .io_in_shift(PE_Array_23_7_io_in_shift),
    .io_out_activate(PE_Array_23_7_io_out_activate),
    .io_out_weight(PE_Array_23_7_io_out_weight),
    .io_out_psum(PE_Array_23_7_io_out_psum)
  );
  basic_PE PE_Array_23_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_8_clock),
    .reset(PE_Array_23_8_reset),
    .io_in_activate(PE_Array_23_8_io_in_activate),
    .io_in_weight(PE_Array_23_8_io_in_weight),
    .io_in_psum(PE_Array_23_8_io_in_psum),
    .io_in_flow(PE_Array_23_8_io_in_flow),
    .io_in_shift(PE_Array_23_8_io_in_shift),
    .io_out_activate(PE_Array_23_8_io_out_activate),
    .io_out_weight(PE_Array_23_8_io_out_weight),
    .io_out_psum(PE_Array_23_8_io_out_psum)
  );
  basic_PE PE_Array_23_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_9_clock),
    .reset(PE_Array_23_9_reset),
    .io_in_activate(PE_Array_23_9_io_in_activate),
    .io_in_weight(PE_Array_23_9_io_in_weight),
    .io_in_psum(PE_Array_23_9_io_in_psum),
    .io_in_flow(PE_Array_23_9_io_in_flow),
    .io_in_shift(PE_Array_23_9_io_in_shift),
    .io_out_activate(PE_Array_23_9_io_out_activate),
    .io_out_weight(PE_Array_23_9_io_out_weight),
    .io_out_psum(PE_Array_23_9_io_out_psum)
  );
  basic_PE PE_Array_23_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_10_clock),
    .reset(PE_Array_23_10_reset),
    .io_in_activate(PE_Array_23_10_io_in_activate),
    .io_in_weight(PE_Array_23_10_io_in_weight),
    .io_in_psum(PE_Array_23_10_io_in_psum),
    .io_in_flow(PE_Array_23_10_io_in_flow),
    .io_in_shift(PE_Array_23_10_io_in_shift),
    .io_out_activate(PE_Array_23_10_io_out_activate),
    .io_out_weight(PE_Array_23_10_io_out_weight),
    .io_out_psum(PE_Array_23_10_io_out_psum)
  );
  basic_PE PE_Array_23_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_11_clock),
    .reset(PE_Array_23_11_reset),
    .io_in_activate(PE_Array_23_11_io_in_activate),
    .io_in_weight(PE_Array_23_11_io_in_weight),
    .io_in_psum(PE_Array_23_11_io_in_psum),
    .io_in_flow(PE_Array_23_11_io_in_flow),
    .io_in_shift(PE_Array_23_11_io_in_shift),
    .io_out_activate(PE_Array_23_11_io_out_activate),
    .io_out_weight(PE_Array_23_11_io_out_weight),
    .io_out_psum(PE_Array_23_11_io_out_psum)
  );
  basic_PE PE_Array_23_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_12_clock),
    .reset(PE_Array_23_12_reset),
    .io_in_activate(PE_Array_23_12_io_in_activate),
    .io_in_weight(PE_Array_23_12_io_in_weight),
    .io_in_psum(PE_Array_23_12_io_in_psum),
    .io_in_flow(PE_Array_23_12_io_in_flow),
    .io_in_shift(PE_Array_23_12_io_in_shift),
    .io_out_activate(PE_Array_23_12_io_out_activate),
    .io_out_weight(PE_Array_23_12_io_out_weight),
    .io_out_psum(PE_Array_23_12_io_out_psum)
  );
  basic_PE PE_Array_23_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_13_clock),
    .reset(PE_Array_23_13_reset),
    .io_in_activate(PE_Array_23_13_io_in_activate),
    .io_in_weight(PE_Array_23_13_io_in_weight),
    .io_in_psum(PE_Array_23_13_io_in_psum),
    .io_in_flow(PE_Array_23_13_io_in_flow),
    .io_in_shift(PE_Array_23_13_io_in_shift),
    .io_out_activate(PE_Array_23_13_io_out_activate),
    .io_out_weight(PE_Array_23_13_io_out_weight),
    .io_out_psum(PE_Array_23_13_io_out_psum)
  );
  basic_PE PE_Array_23_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_14_clock),
    .reset(PE_Array_23_14_reset),
    .io_in_activate(PE_Array_23_14_io_in_activate),
    .io_in_weight(PE_Array_23_14_io_in_weight),
    .io_in_psum(PE_Array_23_14_io_in_psum),
    .io_in_flow(PE_Array_23_14_io_in_flow),
    .io_in_shift(PE_Array_23_14_io_in_shift),
    .io_out_activate(PE_Array_23_14_io_out_activate),
    .io_out_weight(PE_Array_23_14_io_out_weight),
    .io_out_psum(PE_Array_23_14_io_out_psum)
  );
  basic_PE PE_Array_23_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_15_clock),
    .reset(PE_Array_23_15_reset),
    .io_in_activate(PE_Array_23_15_io_in_activate),
    .io_in_weight(PE_Array_23_15_io_in_weight),
    .io_in_psum(PE_Array_23_15_io_in_psum),
    .io_in_flow(PE_Array_23_15_io_in_flow),
    .io_in_shift(PE_Array_23_15_io_in_shift),
    .io_out_activate(PE_Array_23_15_io_out_activate),
    .io_out_weight(PE_Array_23_15_io_out_weight),
    .io_out_psum(PE_Array_23_15_io_out_psum)
  );
  basic_PE PE_Array_23_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_16_clock),
    .reset(PE_Array_23_16_reset),
    .io_in_activate(PE_Array_23_16_io_in_activate),
    .io_in_weight(PE_Array_23_16_io_in_weight),
    .io_in_psum(PE_Array_23_16_io_in_psum),
    .io_in_flow(PE_Array_23_16_io_in_flow),
    .io_in_shift(PE_Array_23_16_io_in_shift),
    .io_out_activate(PE_Array_23_16_io_out_activate),
    .io_out_weight(PE_Array_23_16_io_out_weight),
    .io_out_psum(PE_Array_23_16_io_out_psum)
  );
  basic_PE PE_Array_23_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_17_clock),
    .reset(PE_Array_23_17_reset),
    .io_in_activate(PE_Array_23_17_io_in_activate),
    .io_in_weight(PE_Array_23_17_io_in_weight),
    .io_in_psum(PE_Array_23_17_io_in_psum),
    .io_in_flow(PE_Array_23_17_io_in_flow),
    .io_in_shift(PE_Array_23_17_io_in_shift),
    .io_out_activate(PE_Array_23_17_io_out_activate),
    .io_out_weight(PE_Array_23_17_io_out_weight),
    .io_out_psum(PE_Array_23_17_io_out_psum)
  );
  basic_PE PE_Array_23_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_18_clock),
    .reset(PE_Array_23_18_reset),
    .io_in_activate(PE_Array_23_18_io_in_activate),
    .io_in_weight(PE_Array_23_18_io_in_weight),
    .io_in_psum(PE_Array_23_18_io_in_psum),
    .io_in_flow(PE_Array_23_18_io_in_flow),
    .io_in_shift(PE_Array_23_18_io_in_shift),
    .io_out_activate(PE_Array_23_18_io_out_activate),
    .io_out_weight(PE_Array_23_18_io_out_weight),
    .io_out_psum(PE_Array_23_18_io_out_psum)
  );
  basic_PE PE_Array_23_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_19_clock),
    .reset(PE_Array_23_19_reset),
    .io_in_activate(PE_Array_23_19_io_in_activate),
    .io_in_weight(PE_Array_23_19_io_in_weight),
    .io_in_psum(PE_Array_23_19_io_in_psum),
    .io_in_flow(PE_Array_23_19_io_in_flow),
    .io_in_shift(PE_Array_23_19_io_in_shift),
    .io_out_activate(PE_Array_23_19_io_out_activate),
    .io_out_weight(PE_Array_23_19_io_out_weight),
    .io_out_psum(PE_Array_23_19_io_out_psum)
  );
  basic_PE PE_Array_23_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_20_clock),
    .reset(PE_Array_23_20_reset),
    .io_in_activate(PE_Array_23_20_io_in_activate),
    .io_in_weight(PE_Array_23_20_io_in_weight),
    .io_in_psum(PE_Array_23_20_io_in_psum),
    .io_in_flow(PE_Array_23_20_io_in_flow),
    .io_in_shift(PE_Array_23_20_io_in_shift),
    .io_out_activate(PE_Array_23_20_io_out_activate),
    .io_out_weight(PE_Array_23_20_io_out_weight),
    .io_out_psum(PE_Array_23_20_io_out_psum)
  );
  basic_PE PE_Array_23_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_21_clock),
    .reset(PE_Array_23_21_reset),
    .io_in_activate(PE_Array_23_21_io_in_activate),
    .io_in_weight(PE_Array_23_21_io_in_weight),
    .io_in_psum(PE_Array_23_21_io_in_psum),
    .io_in_flow(PE_Array_23_21_io_in_flow),
    .io_in_shift(PE_Array_23_21_io_in_shift),
    .io_out_activate(PE_Array_23_21_io_out_activate),
    .io_out_weight(PE_Array_23_21_io_out_weight),
    .io_out_psum(PE_Array_23_21_io_out_psum)
  );
  basic_PE PE_Array_23_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_22_clock),
    .reset(PE_Array_23_22_reset),
    .io_in_activate(PE_Array_23_22_io_in_activate),
    .io_in_weight(PE_Array_23_22_io_in_weight),
    .io_in_psum(PE_Array_23_22_io_in_psum),
    .io_in_flow(PE_Array_23_22_io_in_flow),
    .io_in_shift(PE_Array_23_22_io_in_shift),
    .io_out_activate(PE_Array_23_22_io_out_activate),
    .io_out_weight(PE_Array_23_22_io_out_weight),
    .io_out_psum(PE_Array_23_22_io_out_psum)
  );
  basic_PE PE_Array_23_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_23_clock),
    .reset(PE_Array_23_23_reset),
    .io_in_activate(PE_Array_23_23_io_in_activate),
    .io_in_weight(PE_Array_23_23_io_in_weight),
    .io_in_psum(PE_Array_23_23_io_in_psum),
    .io_in_flow(PE_Array_23_23_io_in_flow),
    .io_in_shift(PE_Array_23_23_io_in_shift),
    .io_out_activate(PE_Array_23_23_io_out_activate),
    .io_out_weight(PE_Array_23_23_io_out_weight),
    .io_out_psum(PE_Array_23_23_io_out_psum)
  );
  basic_PE PE_Array_23_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_24_clock),
    .reset(PE_Array_23_24_reset),
    .io_in_activate(PE_Array_23_24_io_in_activate),
    .io_in_weight(PE_Array_23_24_io_in_weight),
    .io_in_psum(PE_Array_23_24_io_in_psum),
    .io_in_flow(PE_Array_23_24_io_in_flow),
    .io_in_shift(PE_Array_23_24_io_in_shift),
    .io_out_activate(PE_Array_23_24_io_out_activate),
    .io_out_weight(PE_Array_23_24_io_out_weight),
    .io_out_psum(PE_Array_23_24_io_out_psum)
  );
  basic_PE PE_Array_23_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_25_clock),
    .reset(PE_Array_23_25_reset),
    .io_in_activate(PE_Array_23_25_io_in_activate),
    .io_in_weight(PE_Array_23_25_io_in_weight),
    .io_in_psum(PE_Array_23_25_io_in_psum),
    .io_in_flow(PE_Array_23_25_io_in_flow),
    .io_in_shift(PE_Array_23_25_io_in_shift),
    .io_out_activate(PE_Array_23_25_io_out_activate),
    .io_out_weight(PE_Array_23_25_io_out_weight),
    .io_out_psum(PE_Array_23_25_io_out_psum)
  );
  basic_PE PE_Array_23_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_26_clock),
    .reset(PE_Array_23_26_reset),
    .io_in_activate(PE_Array_23_26_io_in_activate),
    .io_in_weight(PE_Array_23_26_io_in_weight),
    .io_in_psum(PE_Array_23_26_io_in_psum),
    .io_in_flow(PE_Array_23_26_io_in_flow),
    .io_in_shift(PE_Array_23_26_io_in_shift),
    .io_out_activate(PE_Array_23_26_io_out_activate),
    .io_out_weight(PE_Array_23_26_io_out_weight),
    .io_out_psum(PE_Array_23_26_io_out_psum)
  );
  basic_PE PE_Array_23_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_27_clock),
    .reset(PE_Array_23_27_reset),
    .io_in_activate(PE_Array_23_27_io_in_activate),
    .io_in_weight(PE_Array_23_27_io_in_weight),
    .io_in_psum(PE_Array_23_27_io_in_psum),
    .io_in_flow(PE_Array_23_27_io_in_flow),
    .io_in_shift(PE_Array_23_27_io_in_shift),
    .io_out_activate(PE_Array_23_27_io_out_activate),
    .io_out_weight(PE_Array_23_27_io_out_weight),
    .io_out_psum(PE_Array_23_27_io_out_psum)
  );
  basic_PE PE_Array_23_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_28_clock),
    .reset(PE_Array_23_28_reset),
    .io_in_activate(PE_Array_23_28_io_in_activate),
    .io_in_weight(PE_Array_23_28_io_in_weight),
    .io_in_psum(PE_Array_23_28_io_in_psum),
    .io_in_flow(PE_Array_23_28_io_in_flow),
    .io_in_shift(PE_Array_23_28_io_in_shift),
    .io_out_activate(PE_Array_23_28_io_out_activate),
    .io_out_weight(PE_Array_23_28_io_out_weight),
    .io_out_psum(PE_Array_23_28_io_out_psum)
  );
  basic_PE PE_Array_23_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_29_clock),
    .reset(PE_Array_23_29_reset),
    .io_in_activate(PE_Array_23_29_io_in_activate),
    .io_in_weight(PE_Array_23_29_io_in_weight),
    .io_in_psum(PE_Array_23_29_io_in_psum),
    .io_in_flow(PE_Array_23_29_io_in_flow),
    .io_in_shift(PE_Array_23_29_io_in_shift),
    .io_out_activate(PE_Array_23_29_io_out_activate),
    .io_out_weight(PE_Array_23_29_io_out_weight),
    .io_out_psum(PE_Array_23_29_io_out_psum)
  );
  basic_PE PE_Array_23_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_30_clock),
    .reset(PE_Array_23_30_reset),
    .io_in_activate(PE_Array_23_30_io_in_activate),
    .io_in_weight(PE_Array_23_30_io_in_weight),
    .io_in_psum(PE_Array_23_30_io_in_psum),
    .io_in_flow(PE_Array_23_30_io_in_flow),
    .io_in_shift(PE_Array_23_30_io_in_shift),
    .io_out_activate(PE_Array_23_30_io_out_activate),
    .io_out_weight(PE_Array_23_30_io_out_weight),
    .io_out_psum(PE_Array_23_30_io_out_psum)
  );
  basic_PE PE_Array_23_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_23_31_clock),
    .reset(PE_Array_23_31_reset),
    .io_in_activate(PE_Array_23_31_io_in_activate),
    .io_in_weight(PE_Array_23_31_io_in_weight),
    .io_in_psum(PE_Array_23_31_io_in_psum),
    .io_in_flow(PE_Array_23_31_io_in_flow),
    .io_in_shift(PE_Array_23_31_io_in_shift),
    .io_out_activate(PE_Array_23_31_io_out_activate),
    .io_out_weight(PE_Array_23_31_io_out_weight),
    .io_out_psum(PE_Array_23_31_io_out_psum)
  );
  basic_PE PE_Array_24_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_0_clock),
    .reset(PE_Array_24_0_reset),
    .io_in_activate(PE_Array_24_0_io_in_activate),
    .io_in_weight(PE_Array_24_0_io_in_weight),
    .io_in_psum(PE_Array_24_0_io_in_psum),
    .io_in_flow(PE_Array_24_0_io_in_flow),
    .io_in_shift(PE_Array_24_0_io_in_shift),
    .io_out_activate(PE_Array_24_0_io_out_activate),
    .io_out_weight(PE_Array_24_0_io_out_weight),
    .io_out_psum(PE_Array_24_0_io_out_psum)
  );
  basic_PE PE_Array_24_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_1_clock),
    .reset(PE_Array_24_1_reset),
    .io_in_activate(PE_Array_24_1_io_in_activate),
    .io_in_weight(PE_Array_24_1_io_in_weight),
    .io_in_psum(PE_Array_24_1_io_in_psum),
    .io_in_flow(PE_Array_24_1_io_in_flow),
    .io_in_shift(PE_Array_24_1_io_in_shift),
    .io_out_activate(PE_Array_24_1_io_out_activate),
    .io_out_weight(PE_Array_24_1_io_out_weight),
    .io_out_psum(PE_Array_24_1_io_out_psum)
  );
  basic_PE PE_Array_24_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_2_clock),
    .reset(PE_Array_24_2_reset),
    .io_in_activate(PE_Array_24_2_io_in_activate),
    .io_in_weight(PE_Array_24_2_io_in_weight),
    .io_in_psum(PE_Array_24_2_io_in_psum),
    .io_in_flow(PE_Array_24_2_io_in_flow),
    .io_in_shift(PE_Array_24_2_io_in_shift),
    .io_out_activate(PE_Array_24_2_io_out_activate),
    .io_out_weight(PE_Array_24_2_io_out_weight),
    .io_out_psum(PE_Array_24_2_io_out_psum)
  );
  basic_PE PE_Array_24_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_3_clock),
    .reset(PE_Array_24_3_reset),
    .io_in_activate(PE_Array_24_3_io_in_activate),
    .io_in_weight(PE_Array_24_3_io_in_weight),
    .io_in_psum(PE_Array_24_3_io_in_psum),
    .io_in_flow(PE_Array_24_3_io_in_flow),
    .io_in_shift(PE_Array_24_3_io_in_shift),
    .io_out_activate(PE_Array_24_3_io_out_activate),
    .io_out_weight(PE_Array_24_3_io_out_weight),
    .io_out_psum(PE_Array_24_3_io_out_psum)
  );
  basic_PE PE_Array_24_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_4_clock),
    .reset(PE_Array_24_4_reset),
    .io_in_activate(PE_Array_24_4_io_in_activate),
    .io_in_weight(PE_Array_24_4_io_in_weight),
    .io_in_psum(PE_Array_24_4_io_in_psum),
    .io_in_flow(PE_Array_24_4_io_in_flow),
    .io_in_shift(PE_Array_24_4_io_in_shift),
    .io_out_activate(PE_Array_24_4_io_out_activate),
    .io_out_weight(PE_Array_24_4_io_out_weight),
    .io_out_psum(PE_Array_24_4_io_out_psum)
  );
  basic_PE PE_Array_24_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_5_clock),
    .reset(PE_Array_24_5_reset),
    .io_in_activate(PE_Array_24_5_io_in_activate),
    .io_in_weight(PE_Array_24_5_io_in_weight),
    .io_in_psum(PE_Array_24_5_io_in_psum),
    .io_in_flow(PE_Array_24_5_io_in_flow),
    .io_in_shift(PE_Array_24_5_io_in_shift),
    .io_out_activate(PE_Array_24_5_io_out_activate),
    .io_out_weight(PE_Array_24_5_io_out_weight),
    .io_out_psum(PE_Array_24_5_io_out_psum)
  );
  basic_PE PE_Array_24_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_6_clock),
    .reset(PE_Array_24_6_reset),
    .io_in_activate(PE_Array_24_6_io_in_activate),
    .io_in_weight(PE_Array_24_6_io_in_weight),
    .io_in_psum(PE_Array_24_6_io_in_psum),
    .io_in_flow(PE_Array_24_6_io_in_flow),
    .io_in_shift(PE_Array_24_6_io_in_shift),
    .io_out_activate(PE_Array_24_6_io_out_activate),
    .io_out_weight(PE_Array_24_6_io_out_weight),
    .io_out_psum(PE_Array_24_6_io_out_psum)
  );
  basic_PE PE_Array_24_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_7_clock),
    .reset(PE_Array_24_7_reset),
    .io_in_activate(PE_Array_24_7_io_in_activate),
    .io_in_weight(PE_Array_24_7_io_in_weight),
    .io_in_psum(PE_Array_24_7_io_in_psum),
    .io_in_flow(PE_Array_24_7_io_in_flow),
    .io_in_shift(PE_Array_24_7_io_in_shift),
    .io_out_activate(PE_Array_24_7_io_out_activate),
    .io_out_weight(PE_Array_24_7_io_out_weight),
    .io_out_psum(PE_Array_24_7_io_out_psum)
  );
  basic_PE PE_Array_24_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_8_clock),
    .reset(PE_Array_24_8_reset),
    .io_in_activate(PE_Array_24_8_io_in_activate),
    .io_in_weight(PE_Array_24_8_io_in_weight),
    .io_in_psum(PE_Array_24_8_io_in_psum),
    .io_in_flow(PE_Array_24_8_io_in_flow),
    .io_in_shift(PE_Array_24_8_io_in_shift),
    .io_out_activate(PE_Array_24_8_io_out_activate),
    .io_out_weight(PE_Array_24_8_io_out_weight),
    .io_out_psum(PE_Array_24_8_io_out_psum)
  );
  basic_PE PE_Array_24_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_9_clock),
    .reset(PE_Array_24_9_reset),
    .io_in_activate(PE_Array_24_9_io_in_activate),
    .io_in_weight(PE_Array_24_9_io_in_weight),
    .io_in_psum(PE_Array_24_9_io_in_psum),
    .io_in_flow(PE_Array_24_9_io_in_flow),
    .io_in_shift(PE_Array_24_9_io_in_shift),
    .io_out_activate(PE_Array_24_9_io_out_activate),
    .io_out_weight(PE_Array_24_9_io_out_weight),
    .io_out_psum(PE_Array_24_9_io_out_psum)
  );
  basic_PE PE_Array_24_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_10_clock),
    .reset(PE_Array_24_10_reset),
    .io_in_activate(PE_Array_24_10_io_in_activate),
    .io_in_weight(PE_Array_24_10_io_in_weight),
    .io_in_psum(PE_Array_24_10_io_in_psum),
    .io_in_flow(PE_Array_24_10_io_in_flow),
    .io_in_shift(PE_Array_24_10_io_in_shift),
    .io_out_activate(PE_Array_24_10_io_out_activate),
    .io_out_weight(PE_Array_24_10_io_out_weight),
    .io_out_psum(PE_Array_24_10_io_out_psum)
  );
  basic_PE PE_Array_24_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_11_clock),
    .reset(PE_Array_24_11_reset),
    .io_in_activate(PE_Array_24_11_io_in_activate),
    .io_in_weight(PE_Array_24_11_io_in_weight),
    .io_in_psum(PE_Array_24_11_io_in_psum),
    .io_in_flow(PE_Array_24_11_io_in_flow),
    .io_in_shift(PE_Array_24_11_io_in_shift),
    .io_out_activate(PE_Array_24_11_io_out_activate),
    .io_out_weight(PE_Array_24_11_io_out_weight),
    .io_out_psum(PE_Array_24_11_io_out_psum)
  );
  basic_PE PE_Array_24_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_12_clock),
    .reset(PE_Array_24_12_reset),
    .io_in_activate(PE_Array_24_12_io_in_activate),
    .io_in_weight(PE_Array_24_12_io_in_weight),
    .io_in_psum(PE_Array_24_12_io_in_psum),
    .io_in_flow(PE_Array_24_12_io_in_flow),
    .io_in_shift(PE_Array_24_12_io_in_shift),
    .io_out_activate(PE_Array_24_12_io_out_activate),
    .io_out_weight(PE_Array_24_12_io_out_weight),
    .io_out_psum(PE_Array_24_12_io_out_psum)
  );
  basic_PE PE_Array_24_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_13_clock),
    .reset(PE_Array_24_13_reset),
    .io_in_activate(PE_Array_24_13_io_in_activate),
    .io_in_weight(PE_Array_24_13_io_in_weight),
    .io_in_psum(PE_Array_24_13_io_in_psum),
    .io_in_flow(PE_Array_24_13_io_in_flow),
    .io_in_shift(PE_Array_24_13_io_in_shift),
    .io_out_activate(PE_Array_24_13_io_out_activate),
    .io_out_weight(PE_Array_24_13_io_out_weight),
    .io_out_psum(PE_Array_24_13_io_out_psum)
  );
  basic_PE PE_Array_24_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_14_clock),
    .reset(PE_Array_24_14_reset),
    .io_in_activate(PE_Array_24_14_io_in_activate),
    .io_in_weight(PE_Array_24_14_io_in_weight),
    .io_in_psum(PE_Array_24_14_io_in_psum),
    .io_in_flow(PE_Array_24_14_io_in_flow),
    .io_in_shift(PE_Array_24_14_io_in_shift),
    .io_out_activate(PE_Array_24_14_io_out_activate),
    .io_out_weight(PE_Array_24_14_io_out_weight),
    .io_out_psum(PE_Array_24_14_io_out_psum)
  );
  basic_PE PE_Array_24_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_15_clock),
    .reset(PE_Array_24_15_reset),
    .io_in_activate(PE_Array_24_15_io_in_activate),
    .io_in_weight(PE_Array_24_15_io_in_weight),
    .io_in_psum(PE_Array_24_15_io_in_psum),
    .io_in_flow(PE_Array_24_15_io_in_flow),
    .io_in_shift(PE_Array_24_15_io_in_shift),
    .io_out_activate(PE_Array_24_15_io_out_activate),
    .io_out_weight(PE_Array_24_15_io_out_weight),
    .io_out_psum(PE_Array_24_15_io_out_psum)
  );
  basic_PE PE_Array_24_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_16_clock),
    .reset(PE_Array_24_16_reset),
    .io_in_activate(PE_Array_24_16_io_in_activate),
    .io_in_weight(PE_Array_24_16_io_in_weight),
    .io_in_psum(PE_Array_24_16_io_in_psum),
    .io_in_flow(PE_Array_24_16_io_in_flow),
    .io_in_shift(PE_Array_24_16_io_in_shift),
    .io_out_activate(PE_Array_24_16_io_out_activate),
    .io_out_weight(PE_Array_24_16_io_out_weight),
    .io_out_psum(PE_Array_24_16_io_out_psum)
  );
  basic_PE PE_Array_24_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_17_clock),
    .reset(PE_Array_24_17_reset),
    .io_in_activate(PE_Array_24_17_io_in_activate),
    .io_in_weight(PE_Array_24_17_io_in_weight),
    .io_in_psum(PE_Array_24_17_io_in_psum),
    .io_in_flow(PE_Array_24_17_io_in_flow),
    .io_in_shift(PE_Array_24_17_io_in_shift),
    .io_out_activate(PE_Array_24_17_io_out_activate),
    .io_out_weight(PE_Array_24_17_io_out_weight),
    .io_out_psum(PE_Array_24_17_io_out_psum)
  );
  basic_PE PE_Array_24_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_18_clock),
    .reset(PE_Array_24_18_reset),
    .io_in_activate(PE_Array_24_18_io_in_activate),
    .io_in_weight(PE_Array_24_18_io_in_weight),
    .io_in_psum(PE_Array_24_18_io_in_psum),
    .io_in_flow(PE_Array_24_18_io_in_flow),
    .io_in_shift(PE_Array_24_18_io_in_shift),
    .io_out_activate(PE_Array_24_18_io_out_activate),
    .io_out_weight(PE_Array_24_18_io_out_weight),
    .io_out_psum(PE_Array_24_18_io_out_psum)
  );
  basic_PE PE_Array_24_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_19_clock),
    .reset(PE_Array_24_19_reset),
    .io_in_activate(PE_Array_24_19_io_in_activate),
    .io_in_weight(PE_Array_24_19_io_in_weight),
    .io_in_psum(PE_Array_24_19_io_in_psum),
    .io_in_flow(PE_Array_24_19_io_in_flow),
    .io_in_shift(PE_Array_24_19_io_in_shift),
    .io_out_activate(PE_Array_24_19_io_out_activate),
    .io_out_weight(PE_Array_24_19_io_out_weight),
    .io_out_psum(PE_Array_24_19_io_out_psum)
  );
  basic_PE PE_Array_24_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_20_clock),
    .reset(PE_Array_24_20_reset),
    .io_in_activate(PE_Array_24_20_io_in_activate),
    .io_in_weight(PE_Array_24_20_io_in_weight),
    .io_in_psum(PE_Array_24_20_io_in_psum),
    .io_in_flow(PE_Array_24_20_io_in_flow),
    .io_in_shift(PE_Array_24_20_io_in_shift),
    .io_out_activate(PE_Array_24_20_io_out_activate),
    .io_out_weight(PE_Array_24_20_io_out_weight),
    .io_out_psum(PE_Array_24_20_io_out_psum)
  );
  basic_PE PE_Array_24_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_21_clock),
    .reset(PE_Array_24_21_reset),
    .io_in_activate(PE_Array_24_21_io_in_activate),
    .io_in_weight(PE_Array_24_21_io_in_weight),
    .io_in_psum(PE_Array_24_21_io_in_psum),
    .io_in_flow(PE_Array_24_21_io_in_flow),
    .io_in_shift(PE_Array_24_21_io_in_shift),
    .io_out_activate(PE_Array_24_21_io_out_activate),
    .io_out_weight(PE_Array_24_21_io_out_weight),
    .io_out_psum(PE_Array_24_21_io_out_psum)
  );
  basic_PE PE_Array_24_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_22_clock),
    .reset(PE_Array_24_22_reset),
    .io_in_activate(PE_Array_24_22_io_in_activate),
    .io_in_weight(PE_Array_24_22_io_in_weight),
    .io_in_psum(PE_Array_24_22_io_in_psum),
    .io_in_flow(PE_Array_24_22_io_in_flow),
    .io_in_shift(PE_Array_24_22_io_in_shift),
    .io_out_activate(PE_Array_24_22_io_out_activate),
    .io_out_weight(PE_Array_24_22_io_out_weight),
    .io_out_psum(PE_Array_24_22_io_out_psum)
  );
  basic_PE PE_Array_24_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_23_clock),
    .reset(PE_Array_24_23_reset),
    .io_in_activate(PE_Array_24_23_io_in_activate),
    .io_in_weight(PE_Array_24_23_io_in_weight),
    .io_in_psum(PE_Array_24_23_io_in_psum),
    .io_in_flow(PE_Array_24_23_io_in_flow),
    .io_in_shift(PE_Array_24_23_io_in_shift),
    .io_out_activate(PE_Array_24_23_io_out_activate),
    .io_out_weight(PE_Array_24_23_io_out_weight),
    .io_out_psum(PE_Array_24_23_io_out_psum)
  );
  basic_PE PE_Array_24_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_24_clock),
    .reset(PE_Array_24_24_reset),
    .io_in_activate(PE_Array_24_24_io_in_activate),
    .io_in_weight(PE_Array_24_24_io_in_weight),
    .io_in_psum(PE_Array_24_24_io_in_psum),
    .io_in_flow(PE_Array_24_24_io_in_flow),
    .io_in_shift(PE_Array_24_24_io_in_shift),
    .io_out_activate(PE_Array_24_24_io_out_activate),
    .io_out_weight(PE_Array_24_24_io_out_weight),
    .io_out_psum(PE_Array_24_24_io_out_psum)
  );
  basic_PE PE_Array_24_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_25_clock),
    .reset(PE_Array_24_25_reset),
    .io_in_activate(PE_Array_24_25_io_in_activate),
    .io_in_weight(PE_Array_24_25_io_in_weight),
    .io_in_psum(PE_Array_24_25_io_in_psum),
    .io_in_flow(PE_Array_24_25_io_in_flow),
    .io_in_shift(PE_Array_24_25_io_in_shift),
    .io_out_activate(PE_Array_24_25_io_out_activate),
    .io_out_weight(PE_Array_24_25_io_out_weight),
    .io_out_psum(PE_Array_24_25_io_out_psum)
  );
  basic_PE PE_Array_24_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_26_clock),
    .reset(PE_Array_24_26_reset),
    .io_in_activate(PE_Array_24_26_io_in_activate),
    .io_in_weight(PE_Array_24_26_io_in_weight),
    .io_in_psum(PE_Array_24_26_io_in_psum),
    .io_in_flow(PE_Array_24_26_io_in_flow),
    .io_in_shift(PE_Array_24_26_io_in_shift),
    .io_out_activate(PE_Array_24_26_io_out_activate),
    .io_out_weight(PE_Array_24_26_io_out_weight),
    .io_out_psum(PE_Array_24_26_io_out_psum)
  );
  basic_PE PE_Array_24_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_27_clock),
    .reset(PE_Array_24_27_reset),
    .io_in_activate(PE_Array_24_27_io_in_activate),
    .io_in_weight(PE_Array_24_27_io_in_weight),
    .io_in_psum(PE_Array_24_27_io_in_psum),
    .io_in_flow(PE_Array_24_27_io_in_flow),
    .io_in_shift(PE_Array_24_27_io_in_shift),
    .io_out_activate(PE_Array_24_27_io_out_activate),
    .io_out_weight(PE_Array_24_27_io_out_weight),
    .io_out_psum(PE_Array_24_27_io_out_psum)
  );
  basic_PE PE_Array_24_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_28_clock),
    .reset(PE_Array_24_28_reset),
    .io_in_activate(PE_Array_24_28_io_in_activate),
    .io_in_weight(PE_Array_24_28_io_in_weight),
    .io_in_psum(PE_Array_24_28_io_in_psum),
    .io_in_flow(PE_Array_24_28_io_in_flow),
    .io_in_shift(PE_Array_24_28_io_in_shift),
    .io_out_activate(PE_Array_24_28_io_out_activate),
    .io_out_weight(PE_Array_24_28_io_out_weight),
    .io_out_psum(PE_Array_24_28_io_out_psum)
  );
  basic_PE PE_Array_24_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_29_clock),
    .reset(PE_Array_24_29_reset),
    .io_in_activate(PE_Array_24_29_io_in_activate),
    .io_in_weight(PE_Array_24_29_io_in_weight),
    .io_in_psum(PE_Array_24_29_io_in_psum),
    .io_in_flow(PE_Array_24_29_io_in_flow),
    .io_in_shift(PE_Array_24_29_io_in_shift),
    .io_out_activate(PE_Array_24_29_io_out_activate),
    .io_out_weight(PE_Array_24_29_io_out_weight),
    .io_out_psum(PE_Array_24_29_io_out_psum)
  );
  basic_PE PE_Array_24_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_30_clock),
    .reset(PE_Array_24_30_reset),
    .io_in_activate(PE_Array_24_30_io_in_activate),
    .io_in_weight(PE_Array_24_30_io_in_weight),
    .io_in_psum(PE_Array_24_30_io_in_psum),
    .io_in_flow(PE_Array_24_30_io_in_flow),
    .io_in_shift(PE_Array_24_30_io_in_shift),
    .io_out_activate(PE_Array_24_30_io_out_activate),
    .io_out_weight(PE_Array_24_30_io_out_weight),
    .io_out_psum(PE_Array_24_30_io_out_psum)
  );
  basic_PE PE_Array_24_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_24_31_clock),
    .reset(PE_Array_24_31_reset),
    .io_in_activate(PE_Array_24_31_io_in_activate),
    .io_in_weight(PE_Array_24_31_io_in_weight),
    .io_in_psum(PE_Array_24_31_io_in_psum),
    .io_in_flow(PE_Array_24_31_io_in_flow),
    .io_in_shift(PE_Array_24_31_io_in_shift),
    .io_out_activate(PE_Array_24_31_io_out_activate),
    .io_out_weight(PE_Array_24_31_io_out_weight),
    .io_out_psum(PE_Array_24_31_io_out_psum)
  );
  basic_PE PE_Array_25_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_0_clock),
    .reset(PE_Array_25_0_reset),
    .io_in_activate(PE_Array_25_0_io_in_activate),
    .io_in_weight(PE_Array_25_0_io_in_weight),
    .io_in_psum(PE_Array_25_0_io_in_psum),
    .io_in_flow(PE_Array_25_0_io_in_flow),
    .io_in_shift(PE_Array_25_0_io_in_shift),
    .io_out_activate(PE_Array_25_0_io_out_activate),
    .io_out_weight(PE_Array_25_0_io_out_weight),
    .io_out_psum(PE_Array_25_0_io_out_psum)
  );
  basic_PE PE_Array_25_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_1_clock),
    .reset(PE_Array_25_1_reset),
    .io_in_activate(PE_Array_25_1_io_in_activate),
    .io_in_weight(PE_Array_25_1_io_in_weight),
    .io_in_psum(PE_Array_25_1_io_in_psum),
    .io_in_flow(PE_Array_25_1_io_in_flow),
    .io_in_shift(PE_Array_25_1_io_in_shift),
    .io_out_activate(PE_Array_25_1_io_out_activate),
    .io_out_weight(PE_Array_25_1_io_out_weight),
    .io_out_psum(PE_Array_25_1_io_out_psum)
  );
  basic_PE PE_Array_25_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_2_clock),
    .reset(PE_Array_25_2_reset),
    .io_in_activate(PE_Array_25_2_io_in_activate),
    .io_in_weight(PE_Array_25_2_io_in_weight),
    .io_in_psum(PE_Array_25_2_io_in_psum),
    .io_in_flow(PE_Array_25_2_io_in_flow),
    .io_in_shift(PE_Array_25_2_io_in_shift),
    .io_out_activate(PE_Array_25_2_io_out_activate),
    .io_out_weight(PE_Array_25_2_io_out_weight),
    .io_out_psum(PE_Array_25_2_io_out_psum)
  );
  basic_PE PE_Array_25_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_3_clock),
    .reset(PE_Array_25_3_reset),
    .io_in_activate(PE_Array_25_3_io_in_activate),
    .io_in_weight(PE_Array_25_3_io_in_weight),
    .io_in_psum(PE_Array_25_3_io_in_psum),
    .io_in_flow(PE_Array_25_3_io_in_flow),
    .io_in_shift(PE_Array_25_3_io_in_shift),
    .io_out_activate(PE_Array_25_3_io_out_activate),
    .io_out_weight(PE_Array_25_3_io_out_weight),
    .io_out_psum(PE_Array_25_3_io_out_psum)
  );
  basic_PE PE_Array_25_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_4_clock),
    .reset(PE_Array_25_4_reset),
    .io_in_activate(PE_Array_25_4_io_in_activate),
    .io_in_weight(PE_Array_25_4_io_in_weight),
    .io_in_psum(PE_Array_25_4_io_in_psum),
    .io_in_flow(PE_Array_25_4_io_in_flow),
    .io_in_shift(PE_Array_25_4_io_in_shift),
    .io_out_activate(PE_Array_25_4_io_out_activate),
    .io_out_weight(PE_Array_25_4_io_out_weight),
    .io_out_psum(PE_Array_25_4_io_out_psum)
  );
  basic_PE PE_Array_25_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_5_clock),
    .reset(PE_Array_25_5_reset),
    .io_in_activate(PE_Array_25_5_io_in_activate),
    .io_in_weight(PE_Array_25_5_io_in_weight),
    .io_in_psum(PE_Array_25_5_io_in_psum),
    .io_in_flow(PE_Array_25_5_io_in_flow),
    .io_in_shift(PE_Array_25_5_io_in_shift),
    .io_out_activate(PE_Array_25_5_io_out_activate),
    .io_out_weight(PE_Array_25_5_io_out_weight),
    .io_out_psum(PE_Array_25_5_io_out_psum)
  );
  basic_PE PE_Array_25_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_6_clock),
    .reset(PE_Array_25_6_reset),
    .io_in_activate(PE_Array_25_6_io_in_activate),
    .io_in_weight(PE_Array_25_6_io_in_weight),
    .io_in_psum(PE_Array_25_6_io_in_psum),
    .io_in_flow(PE_Array_25_6_io_in_flow),
    .io_in_shift(PE_Array_25_6_io_in_shift),
    .io_out_activate(PE_Array_25_6_io_out_activate),
    .io_out_weight(PE_Array_25_6_io_out_weight),
    .io_out_psum(PE_Array_25_6_io_out_psum)
  );
  basic_PE PE_Array_25_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_7_clock),
    .reset(PE_Array_25_7_reset),
    .io_in_activate(PE_Array_25_7_io_in_activate),
    .io_in_weight(PE_Array_25_7_io_in_weight),
    .io_in_psum(PE_Array_25_7_io_in_psum),
    .io_in_flow(PE_Array_25_7_io_in_flow),
    .io_in_shift(PE_Array_25_7_io_in_shift),
    .io_out_activate(PE_Array_25_7_io_out_activate),
    .io_out_weight(PE_Array_25_7_io_out_weight),
    .io_out_psum(PE_Array_25_7_io_out_psum)
  );
  basic_PE PE_Array_25_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_8_clock),
    .reset(PE_Array_25_8_reset),
    .io_in_activate(PE_Array_25_8_io_in_activate),
    .io_in_weight(PE_Array_25_8_io_in_weight),
    .io_in_psum(PE_Array_25_8_io_in_psum),
    .io_in_flow(PE_Array_25_8_io_in_flow),
    .io_in_shift(PE_Array_25_8_io_in_shift),
    .io_out_activate(PE_Array_25_8_io_out_activate),
    .io_out_weight(PE_Array_25_8_io_out_weight),
    .io_out_psum(PE_Array_25_8_io_out_psum)
  );
  basic_PE PE_Array_25_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_9_clock),
    .reset(PE_Array_25_9_reset),
    .io_in_activate(PE_Array_25_9_io_in_activate),
    .io_in_weight(PE_Array_25_9_io_in_weight),
    .io_in_psum(PE_Array_25_9_io_in_psum),
    .io_in_flow(PE_Array_25_9_io_in_flow),
    .io_in_shift(PE_Array_25_9_io_in_shift),
    .io_out_activate(PE_Array_25_9_io_out_activate),
    .io_out_weight(PE_Array_25_9_io_out_weight),
    .io_out_psum(PE_Array_25_9_io_out_psum)
  );
  basic_PE PE_Array_25_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_10_clock),
    .reset(PE_Array_25_10_reset),
    .io_in_activate(PE_Array_25_10_io_in_activate),
    .io_in_weight(PE_Array_25_10_io_in_weight),
    .io_in_psum(PE_Array_25_10_io_in_psum),
    .io_in_flow(PE_Array_25_10_io_in_flow),
    .io_in_shift(PE_Array_25_10_io_in_shift),
    .io_out_activate(PE_Array_25_10_io_out_activate),
    .io_out_weight(PE_Array_25_10_io_out_weight),
    .io_out_psum(PE_Array_25_10_io_out_psum)
  );
  basic_PE PE_Array_25_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_11_clock),
    .reset(PE_Array_25_11_reset),
    .io_in_activate(PE_Array_25_11_io_in_activate),
    .io_in_weight(PE_Array_25_11_io_in_weight),
    .io_in_psum(PE_Array_25_11_io_in_psum),
    .io_in_flow(PE_Array_25_11_io_in_flow),
    .io_in_shift(PE_Array_25_11_io_in_shift),
    .io_out_activate(PE_Array_25_11_io_out_activate),
    .io_out_weight(PE_Array_25_11_io_out_weight),
    .io_out_psum(PE_Array_25_11_io_out_psum)
  );
  basic_PE PE_Array_25_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_12_clock),
    .reset(PE_Array_25_12_reset),
    .io_in_activate(PE_Array_25_12_io_in_activate),
    .io_in_weight(PE_Array_25_12_io_in_weight),
    .io_in_psum(PE_Array_25_12_io_in_psum),
    .io_in_flow(PE_Array_25_12_io_in_flow),
    .io_in_shift(PE_Array_25_12_io_in_shift),
    .io_out_activate(PE_Array_25_12_io_out_activate),
    .io_out_weight(PE_Array_25_12_io_out_weight),
    .io_out_psum(PE_Array_25_12_io_out_psum)
  );
  basic_PE PE_Array_25_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_13_clock),
    .reset(PE_Array_25_13_reset),
    .io_in_activate(PE_Array_25_13_io_in_activate),
    .io_in_weight(PE_Array_25_13_io_in_weight),
    .io_in_psum(PE_Array_25_13_io_in_psum),
    .io_in_flow(PE_Array_25_13_io_in_flow),
    .io_in_shift(PE_Array_25_13_io_in_shift),
    .io_out_activate(PE_Array_25_13_io_out_activate),
    .io_out_weight(PE_Array_25_13_io_out_weight),
    .io_out_psum(PE_Array_25_13_io_out_psum)
  );
  basic_PE PE_Array_25_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_14_clock),
    .reset(PE_Array_25_14_reset),
    .io_in_activate(PE_Array_25_14_io_in_activate),
    .io_in_weight(PE_Array_25_14_io_in_weight),
    .io_in_psum(PE_Array_25_14_io_in_psum),
    .io_in_flow(PE_Array_25_14_io_in_flow),
    .io_in_shift(PE_Array_25_14_io_in_shift),
    .io_out_activate(PE_Array_25_14_io_out_activate),
    .io_out_weight(PE_Array_25_14_io_out_weight),
    .io_out_psum(PE_Array_25_14_io_out_psum)
  );
  basic_PE PE_Array_25_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_15_clock),
    .reset(PE_Array_25_15_reset),
    .io_in_activate(PE_Array_25_15_io_in_activate),
    .io_in_weight(PE_Array_25_15_io_in_weight),
    .io_in_psum(PE_Array_25_15_io_in_psum),
    .io_in_flow(PE_Array_25_15_io_in_flow),
    .io_in_shift(PE_Array_25_15_io_in_shift),
    .io_out_activate(PE_Array_25_15_io_out_activate),
    .io_out_weight(PE_Array_25_15_io_out_weight),
    .io_out_psum(PE_Array_25_15_io_out_psum)
  );
  basic_PE PE_Array_25_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_16_clock),
    .reset(PE_Array_25_16_reset),
    .io_in_activate(PE_Array_25_16_io_in_activate),
    .io_in_weight(PE_Array_25_16_io_in_weight),
    .io_in_psum(PE_Array_25_16_io_in_psum),
    .io_in_flow(PE_Array_25_16_io_in_flow),
    .io_in_shift(PE_Array_25_16_io_in_shift),
    .io_out_activate(PE_Array_25_16_io_out_activate),
    .io_out_weight(PE_Array_25_16_io_out_weight),
    .io_out_psum(PE_Array_25_16_io_out_psum)
  );
  basic_PE PE_Array_25_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_17_clock),
    .reset(PE_Array_25_17_reset),
    .io_in_activate(PE_Array_25_17_io_in_activate),
    .io_in_weight(PE_Array_25_17_io_in_weight),
    .io_in_psum(PE_Array_25_17_io_in_psum),
    .io_in_flow(PE_Array_25_17_io_in_flow),
    .io_in_shift(PE_Array_25_17_io_in_shift),
    .io_out_activate(PE_Array_25_17_io_out_activate),
    .io_out_weight(PE_Array_25_17_io_out_weight),
    .io_out_psum(PE_Array_25_17_io_out_psum)
  );
  basic_PE PE_Array_25_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_18_clock),
    .reset(PE_Array_25_18_reset),
    .io_in_activate(PE_Array_25_18_io_in_activate),
    .io_in_weight(PE_Array_25_18_io_in_weight),
    .io_in_psum(PE_Array_25_18_io_in_psum),
    .io_in_flow(PE_Array_25_18_io_in_flow),
    .io_in_shift(PE_Array_25_18_io_in_shift),
    .io_out_activate(PE_Array_25_18_io_out_activate),
    .io_out_weight(PE_Array_25_18_io_out_weight),
    .io_out_psum(PE_Array_25_18_io_out_psum)
  );
  basic_PE PE_Array_25_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_19_clock),
    .reset(PE_Array_25_19_reset),
    .io_in_activate(PE_Array_25_19_io_in_activate),
    .io_in_weight(PE_Array_25_19_io_in_weight),
    .io_in_psum(PE_Array_25_19_io_in_psum),
    .io_in_flow(PE_Array_25_19_io_in_flow),
    .io_in_shift(PE_Array_25_19_io_in_shift),
    .io_out_activate(PE_Array_25_19_io_out_activate),
    .io_out_weight(PE_Array_25_19_io_out_weight),
    .io_out_psum(PE_Array_25_19_io_out_psum)
  );
  basic_PE PE_Array_25_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_20_clock),
    .reset(PE_Array_25_20_reset),
    .io_in_activate(PE_Array_25_20_io_in_activate),
    .io_in_weight(PE_Array_25_20_io_in_weight),
    .io_in_psum(PE_Array_25_20_io_in_psum),
    .io_in_flow(PE_Array_25_20_io_in_flow),
    .io_in_shift(PE_Array_25_20_io_in_shift),
    .io_out_activate(PE_Array_25_20_io_out_activate),
    .io_out_weight(PE_Array_25_20_io_out_weight),
    .io_out_psum(PE_Array_25_20_io_out_psum)
  );
  basic_PE PE_Array_25_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_21_clock),
    .reset(PE_Array_25_21_reset),
    .io_in_activate(PE_Array_25_21_io_in_activate),
    .io_in_weight(PE_Array_25_21_io_in_weight),
    .io_in_psum(PE_Array_25_21_io_in_psum),
    .io_in_flow(PE_Array_25_21_io_in_flow),
    .io_in_shift(PE_Array_25_21_io_in_shift),
    .io_out_activate(PE_Array_25_21_io_out_activate),
    .io_out_weight(PE_Array_25_21_io_out_weight),
    .io_out_psum(PE_Array_25_21_io_out_psum)
  );
  basic_PE PE_Array_25_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_22_clock),
    .reset(PE_Array_25_22_reset),
    .io_in_activate(PE_Array_25_22_io_in_activate),
    .io_in_weight(PE_Array_25_22_io_in_weight),
    .io_in_psum(PE_Array_25_22_io_in_psum),
    .io_in_flow(PE_Array_25_22_io_in_flow),
    .io_in_shift(PE_Array_25_22_io_in_shift),
    .io_out_activate(PE_Array_25_22_io_out_activate),
    .io_out_weight(PE_Array_25_22_io_out_weight),
    .io_out_psum(PE_Array_25_22_io_out_psum)
  );
  basic_PE PE_Array_25_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_23_clock),
    .reset(PE_Array_25_23_reset),
    .io_in_activate(PE_Array_25_23_io_in_activate),
    .io_in_weight(PE_Array_25_23_io_in_weight),
    .io_in_psum(PE_Array_25_23_io_in_psum),
    .io_in_flow(PE_Array_25_23_io_in_flow),
    .io_in_shift(PE_Array_25_23_io_in_shift),
    .io_out_activate(PE_Array_25_23_io_out_activate),
    .io_out_weight(PE_Array_25_23_io_out_weight),
    .io_out_psum(PE_Array_25_23_io_out_psum)
  );
  basic_PE PE_Array_25_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_24_clock),
    .reset(PE_Array_25_24_reset),
    .io_in_activate(PE_Array_25_24_io_in_activate),
    .io_in_weight(PE_Array_25_24_io_in_weight),
    .io_in_psum(PE_Array_25_24_io_in_psum),
    .io_in_flow(PE_Array_25_24_io_in_flow),
    .io_in_shift(PE_Array_25_24_io_in_shift),
    .io_out_activate(PE_Array_25_24_io_out_activate),
    .io_out_weight(PE_Array_25_24_io_out_weight),
    .io_out_psum(PE_Array_25_24_io_out_psum)
  );
  basic_PE PE_Array_25_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_25_clock),
    .reset(PE_Array_25_25_reset),
    .io_in_activate(PE_Array_25_25_io_in_activate),
    .io_in_weight(PE_Array_25_25_io_in_weight),
    .io_in_psum(PE_Array_25_25_io_in_psum),
    .io_in_flow(PE_Array_25_25_io_in_flow),
    .io_in_shift(PE_Array_25_25_io_in_shift),
    .io_out_activate(PE_Array_25_25_io_out_activate),
    .io_out_weight(PE_Array_25_25_io_out_weight),
    .io_out_psum(PE_Array_25_25_io_out_psum)
  );
  basic_PE PE_Array_25_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_26_clock),
    .reset(PE_Array_25_26_reset),
    .io_in_activate(PE_Array_25_26_io_in_activate),
    .io_in_weight(PE_Array_25_26_io_in_weight),
    .io_in_psum(PE_Array_25_26_io_in_psum),
    .io_in_flow(PE_Array_25_26_io_in_flow),
    .io_in_shift(PE_Array_25_26_io_in_shift),
    .io_out_activate(PE_Array_25_26_io_out_activate),
    .io_out_weight(PE_Array_25_26_io_out_weight),
    .io_out_psum(PE_Array_25_26_io_out_psum)
  );
  basic_PE PE_Array_25_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_27_clock),
    .reset(PE_Array_25_27_reset),
    .io_in_activate(PE_Array_25_27_io_in_activate),
    .io_in_weight(PE_Array_25_27_io_in_weight),
    .io_in_psum(PE_Array_25_27_io_in_psum),
    .io_in_flow(PE_Array_25_27_io_in_flow),
    .io_in_shift(PE_Array_25_27_io_in_shift),
    .io_out_activate(PE_Array_25_27_io_out_activate),
    .io_out_weight(PE_Array_25_27_io_out_weight),
    .io_out_psum(PE_Array_25_27_io_out_psum)
  );
  basic_PE PE_Array_25_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_28_clock),
    .reset(PE_Array_25_28_reset),
    .io_in_activate(PE_Array_25_28_io_in_activate),
    .io_in_weight(PE_Array_25_28_io_in_weight),
    .io_in_psum(PE_Array_25_28_io_in_psum),
    .io_in_flow(PE_Array_25_28_io_in_flow),
    .io_in_shift(PE_Array_25_28_io_in_shift),
    .io_out_activate(PE_Array_25_28_io_out_activate),
    .io_out_weight(PE_Array_25_28_io_out_weight),
    .io_out_psum(PE_Array_25_28_io_out_psum)
  );
  basic_PE PE_Array_25_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_29_clock),
    .reset(PE_Array_25_29_reset),
    .io_in_activate(PE_Array_25_29_io_in_activate),
    .io_in_weight(PE_Array_25_29_io_in_weight),
    .io_in_psum(PE_Array_25_29_io_in_psum),
    .io_in_flow(PE_Array_25_29_io_in_flow),
    .io_in_shift(PE_Array_25_29_io_in_shift),
    .io_out_activate(PE_Array_25_29_io_out_activate),
    .io_out_weight(PE_Array_25_29_io_out_weight),
    .io_out_psum(PE_Array_25_29_io_out_psum)
  );
  basic_PE PE_Array_25_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_30_clock),
    .reset(PE_Array_25_30_reset),
    .io_in_activate(PE_Array_25_30_io_in_activate),
    .io_in_weight(PE_Array_25_30_io_in_weight),
    .io_in_psum(PE_Array_25_30_io_in_psum),
    .io_in_flow(PE_Array_25_30_io_in_flow),
    .io_in_shift(PE_Array_25_30_io_in_shift),
    .io_out_activate(PE_Array_25_30_io_out_activate),
    .io_out_weight(PE_Array_25_30_io_out_weight),
    .io_out_psum(PE_Array_25_30_io_out_psum)
  );
  basic_PE PE_Array_25_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_25_31_clock),
    .reset(PE_Array_25_31_reset),
    .io_in_activate(PE_Array_25_31_io_in_activate),
    .io_in_weight(PE_Array_25_31_io_in_weight),
    .io_in_psum(PE_Array_25_31_io_in_psum),
    .io_in_flow(PE_Array_25_31_io_in_flow),
    .io_in_shift(PE_Array_25_31_io_in_shift),
    .io_out_activate(PE_Array_25_31_io_out_activate),
    .io_out_weight(PE_Array_25_31_io_out_weight),
    .io_out_psum(PE_Array_25_31_io_out_psum)
  );
  basic_PE PE_Array_26_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_0_clock),
    .reset(PE_Array_26_0_reset),
    .io_in_activate(PE_Array_26_0_io_in_activate),
    .io_in_weight(PE_Array_26_0_io_in_weight),
    .io_in_psum(PE_Array_26_0_io_in_psum),
    .io_in_flow(PE_Array_26_0_io_in_flow),
    .io_in_shift(PE_Array_26_0_io_in_shift),
    .io_out_activate(PE_Array_26_0_io_out_activate),
    .io_out_weight(PE_Array_26_0_io_out_weight),
    .io_out_psum(PE_Array_26_0_io_out_psum)
  );
  basic_PE PE_Array_26_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_1_clock),
    .reset(PE_Array_26_1_reset),
    .io_in_activate(PE_Array_26_1_io_in_activate),
    .io_in_weight(PE_Array_26_1_io_in_weight),
    .io_in_psum(PE_Array_26_1_io_in_psum),
    .io_in_flow(PE_Array_26_1_io_in_flow),
    .io_in_shift(PE_Array_26_1_io_in_shift),
    .io_out_activate(PE_Array_26_1_io_out_activate),
    .io_out_weight(PE_Array_26_1_io_out_weight),
    .io_out_psum(PE_Array_26_1_io_out_psum)
  );
  basic_PE PE_Array_26_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_2_clock),
    .reset(PE_Array_26_2_reset),
    .io_in_activate(PE_Array_26_2_io_in_activate),
    .io_in_weight(PE_Array_26_2_io_in_weight),
    .io_in_psum(PE_Array_26_2_io_in_psum),
    .io_in_flow(PE_Array_26_2_io_in_flow),
    .io_in_shift(PE_Array_26_2_io_in_shift),
    .io_out_activate(PE_Array_26_2_io_out_activate),
    .io_out_weight(PE_Array_26_2_io_out_weight),
    .io_out_psum(PE_Array_26_2_io_out_psum)
  );
  basic_PE PE_Array_26_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_3_clock),
    .reset(PE_Array_26_3_reset),
    .io_in_activate(PE_Array_26_3_io_in_activate),
    .io_in_weight(PE_Array_26_3_io_in_weight),
    .io_in_psum(PE_Array_26_3_io_in_psum),
    .io_in_flow(PE_Array_26_3_io_in_flow),
    .io_in_shift(PE_Array_26_3_io_in_shift),
    .io_out_activate(PE_Array_26_3_io_out_activate),
    .io_out_weight(PE_Array_26_3_io_out_weight),
    .io_out_psum(PE_Array_26_3_io_out_psum)
  );
  basic_PE PE_Array_26_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_4_clock),
    .reset(PE_Array_26_4_reset),
    .io_in_activate(PE_Array_26_4_io_in_activate),
    .io_in_weight(PE_Array_26_4_io_in_weight),
    .io_in_psum(PE_Array_26_4_io_in_psum),
    .io_in_flow(PE_Array_26_4_io_in_flow),
    .io_in_shift(PE_Array_26_4_io_in_shift),
    .io_out_activate(PE_Array_26_4_io_out_activate),
    .io_out_weight(PE_Array_26_4_io_out_weight),
    .io_out_psum(PE_Array_26_4_io_out_psum)
  );
  basic_PE PE_Array_26_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_5_clock),
    .reset(PE_Array_26_5_reset),
    .io_in_activate(PE_Array_26_5_io_in_activate),
    .io_in_weight(PE_Array_26_5_io_in_weight),
    .io_in_psum(PE_Array_26_5_io_in_psum),
    .io_in_flow(PE_Array_26_5_io_in_flow),
    .io_in_shift(PE_Array_26_5_io_in_shift),
    .io_out_activate(PE_Array_26_5_io_out_activate),
    .io_out_weight(PE_Array_26_5_io_out_weight),
    .io_out_psum(PE_Array_26_5_io_out_psum)
  );
  basic_PE PE_Array_26_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_6_clock),
    .reset(PE_Array_26_6_reset),
    .io_in_activate(PE_Array_26_6_io_in_activate),
    .io_in_weight(PE_Array_26_6_io_in_weight),
    .io_in_psum(PE_Array_26_6_io_in_psum),
    .io_in_flow(PE_Array_26_6_io_in_flow),
    .io_in_shift(PE_Array_26_6_io_in_shift),
    .io_out_activate(PE_Array_26_6_io_out_activate),
    .io_out_weight(PE_Array_26_6_io_out_weight),
    .io_out_psum(PE_Array_26_6_io_out_psum)
  );
  basic_PE PE_Array_26_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_7_clock),
    .reset(PE_Array_26_7_reset),
    .io_in_activate(PE_Array_26_7_io_in_activate),
    .io_in_weight(PE_Array_26_7_io_in_weight),
    .io_in_psum(PE_Array_26_7_io_in_psum),
    .io_in_flow(PE_Array_26_7_io_in_flow),
    .io_in_shift(PE_Array_26_7_io_in_shift),
    .io_out_activate(PE_Array_26_7_io_out_activate),
    .io_out_weight(PE_Array_26_7_io_out_weight),
    .io_out_psum(PE_Array_26_7_io_out_psum)
  );
  basic_PE PE_Array_26_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_8_clock),
    .reset(PE_Array_26_8_reset),
    .io_in_activate(PE_Array_26_8_io_in_activate),
    .io_in_weight(PE_Array_26_8_io_in_weight),
    .io_in_psum(PE_Array_26_8_io_in_psum),
    .io_in_flow(PE_Array_26_8_io_in_flow),
    .io_in_shift(PE_Array_26_8_io_in_shift),
    .io_out_activate(PE_Array_26_8_io_out_activate),
    .io_out_weight(PE_Array_26_8_io_out_weight),
    .io_out_psum(PE_Array_26_8_io_out_psum)
  );
  basic_PE PE_Array_26_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_9_clock),
    .reset(PE_Array_26_9_reset),
    .io_in_activate(PE_Array_26_9_io_in_activate),
    .io_in_weight(PE_Array_26_9_io_in_weight),
    .io_in_psum(PE_Array_26_9_io_in_psum),
    .io_in_flow(PE_Array_26_9_io_in_flow),
    .io_in_shift(PE_Array_26_9_io_in_shift),
    .io_out_activate(PE_Array_26_9_io_out_activate),
    .io_out_weight(PE_Array_26_9_io_out_weight),
    .io_out_psum(PE_Array_26_9_io_out_psum)
  );
  basic_PE PE_Array_26_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_10_clock),
    .reset(PE_Array_26_10_reset),
    .io_in_activate(PE_Array_26_10_io_in_activate),
    .io_in_weight(PE_Array_26_10_io_in_weight),
    .io_in_psum(PE_Array_26_10_io_in_psum),
    .io_in_flow(PE_Array_26_10_io_in_flow),
    .io_in_shift(PE_Array_26_10_io_in_shift),
    .io_out_activate(PE_Array_26_10_io_out_activate),
    .io_out_weight(PE_Array_26_10_io_out_weight),
    .io_out_psum(PE_Array_26_10_io_out_psum)
  );
  basic_PE PE_Array_26_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_11_clock),
    .reset(PE_Array_26_11_reset),
    .io_in_activate(PE_Array_26_11_io_in_activate),
    .io_in_weight(PE_Array_26_11_io_in_weight),
    .io_in_psum(PE_Array_26_11_io_in_psum),
    .io_in_flow(PE_Array_26_11_io_in_flow),
    .io_in_shift(PE_Array_26_11_io_in_shift),
    .io_out_activate(PE_Array_26_11_io_out_activate),
    .io_out_weight(PE_Array_26_11_io_out_weight),
    .io_out_psum(PE_Array_26_11_io_out_psum)
  );
  basic_PE PE_Array_26_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_12_clock),
    .reset(PE_Array_26_12_reset),
    .io_in_activate(PE_Array_26_12_io_in_activate),
    .io_in_weight(PE_Array_26_12_io_in_weight),
    .io_in_psum(PE_Array_26_12_io_in_psum),
    .io_in_flow(PE_Array_26_12_io_in_flow),
    .io_in_shift(PE_Array_26_12_io_in_shift),
    .io_out_activate(PE_Array_26_12_io_out_activate),
    .io_out_weight(PE_Array_26_12_io_out_weight),
    .io_out_psum(PE_Array_26_12_io_out_psum)
  );
  basic_PE PE_Array_26_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_13_clock),
    .reset(PE_Array_26_13_reset),
    .io_in_activate(PE_Array_26_13_io_in_activate),
    .io_in_weight(PE_Array_26_13_io_in_weight),
    .io_in_psum(PE_Array_26_13_io_in_psum),
    .io_in_flow(PE_Array_26_13_io_in_flow),
    .io_in_shift(PE_Array_26_13_io_in_shift),
    .io_out_activate(PE_Array_26_13_io_out_activate),
    .io_out_weight(PE_Array_26_13_io_out_weight),
    .io_out_psum(PE_Array_26_13_io_out_psum)
  );
  basic_PE PE_Array_26_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_14_clock),
    .reset(PE_Array_26_14_reset),
    .io_in_activate(PE_Array_26_14_io_in_activate),
    .io_in_weight(PE_Array_26_14_io_in_weight),
    .io_in_psum(PE_Array_26_14_io_in_psum),
    .io_in_flow(PE_Array_26_14_io_in_flow),
    .io_in_shift(PE_Array_26_14_io_in_shift),
    .io_out_activate(PE_Array_26_14_io_out_activate),
    .io_out_weight(PE_Array_26_14_io_out_weight),
    .io_out_psum(PE_Array_26_14_io_out_psum)
  );
  basic_PE PE_Array_26_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_15_clock),
    .reset(PE_Array_26_15_reset),
    .io_in_activate(PE_Array_26_15_io_in_activate),
    .io_in_weight(PE_Array_26_15_io_in_weight),
    .io_in_psum(PE_Array_26_15_io_in_psum),
    .io_in_flow(PE_Array_26_15_io_in_flow),
    .io_in_shift(PE_Array_26_15_io_in_shift),
    .io_out_activate(PE_Array_26_15_io_out_activate),
    .io_out_weight(PE_Array_26_15_io_out_weight),
    .io_out_psum(PE_Array_26_15_io_out_psum)
  );
  basic_PE PE_Array_26_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_16_clock),
    .reset(PE_Array_26_16_reset),
    .io_in_activate(PE_Array_26_16_io_in_activate),
    .io_in_weight(PE_Array_26_16_io_in_weight),
    .io_in_psum(PE_Array_26_16_io_in_psum),
    .io_in_flow(PE_Array_26_16_io_in_flow),
    .io_in_shift(PE_Array_26_16_io_in_shift),
    .io_out_activate(PE_Array_26_16_io_out_activate),
    .io_out_weight(PE_Array_26_16_io_out_weight),
    .io_out_psum(PE_Array_26_16_io_out_psum)
  );
  basic_PE PE_Array_26_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_17_clock),
    .reset(PE_Array_26_17_reset),
    .io_in_activate(PE_Array_26_17_io_in_activate),
    .io_in_weight(PE_Array_26_17_io_in_weight),
    .io_in_psum(PE_Array_26_17_io_in_psum),
    .io_in_flow(PE_Array_26_17_io_in_flow),
    .io_in_shift(PE_Array_26_17_io_in_shift),
    .io_out_activate(PE_Array_26_17_io_out_activate),
    .io_out_weight(PE_Array_26_17_io_out_weight),
    .io_out_psum(PE_Array_26_17_io_out_psum)
  );
  basic_PE PE_Array_26_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_18_clock),
    .reset(PE_Array_26_18_reset),
    .io_in_activate(PE_Array_26_18_io_in_activate),
    .io_in_weight(PE_Array_26_18_io_in_weight),
    .io_in_psum(PE_Array_26_18_io_in_psum),
    .io_in_flow(PE_Array_26_18_io_in_flow),
    .io_in_shift(PE_Array_26_18_io_in_shift),
    .io_out_activate(PE_Array_26_18_io_out_activate),
    .io_out_weight(PE_Array_26_18_io_out_weight),
    .io_out_psum(PE_Array_26_18_io_out_psum)
  );
  basic_PE PE_Array_26_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_19_clock),
    .reset(PE_Array_26_19_reset),
    .io_in_activate(PE_Array_26_19_io_in_activate),
    .io_in_weight(PE_Array_26_19_io_in_weight),
    .io_in_psum(PE_Array_26_19_io_in_psum),
    .io_in_flow(PE_Array_26_19_io_in_flow),
    .io_in_shift(PE_Array_26_19_io_in_shift),
    .io_out_activate(PE_Array_26_19_io_out_activate),
    .io_out_weight(PE_Array_26_19_io_out_weight),
    .io_out_psum(PE_Array_26_19_io_out_psum)
  );
  basic_PE PE_Array_26_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_20_clock),
    .reset(PE_Array_26_20_reset),
    .io_in_activate(PE_Array_26_20_io_in_activate),
    .io_in_weight(PE_Array_26_20_io_in_weight),
    .io_in_psum(PE_Array_26_20_io_in_psum),
    .io_in_flow(PE_Array_26_20_io_in_flow),
    .io_in_shift(PE_Array_26_20_io_in_shift),
    .io_out_activate(PE_Array_26_20_io_out_activate),
    .io_out_weight(PE_Array_26_20_io_out_weight),
    .io_out_psum(PE_Array_26_20_io_out_psum)
  );
  basic_PE PE_Array_26_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_21_clock),
    .reset(PE_Array_26_21_reset),
    .io_in_activate(PE_Array_26_21_io_in_activate),
    .io_in_weight(PE_Array_26_21_io_in_weight),
    .io_in_psum(PE_Array_26_21_io_in_psum),
    .io_in_flow(PE_Array_26_21_io_in_flow),
    .io_in_shift(PE_Array_26_21_io_in_shift),
    .io_out_activate(PE_Array_26_21_io_out_activate),
    .io_out_weight(PE_Array_26_21_io_out_weight),
    .io_out_psum(PE_Array_26_21_io_out_psum)
  );
  basic_PE PE_Array_26_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_22_clock),
    .reset(PE_Array_26_22_reset),
    .io_in_activate(PE_Array_26_22_io_in_activate),
    .io_in_weight(PE_Array_26_22_io_in_weight),
    .io_in_psum(PE_Array_26_22_io_in_psum),
    .io_in_flow(PE_Array_26_22_io_in_flow),
    .io_in_shift(PE_Array_26_22_io_in_shift),
    .io_out_activate(PE_Array_26_22_io_out_activate),
    .io_out_weight(PE_Array_26_22_io_out_weight),
    .io_out_psum(PE_Array_26_22_io_out_psum)
  );
  basic_PE PE_Array_26_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_23_clock),
    .reset(PE_Array_26_23_reset),
    .io_in_activate(PE_Array_26_23_io_in_activate),
    .io_in_weight(PE_Array_26_23_io_in_weight),
    .io_in_psum(PE_Array_26_23_io_in_psum),
    .io_in_flow(PE_Array_26_23_io_in_flow),
    .io_in_shift(PE_Array_26_23_io_in_shift),
    .io_out_activate(PE_Array_26_23_io_out_activate),
    .io_out_weight(PE_Array_26_23_io_out_weight),
    .io_out_psum(PE_Array_26_23_io_out_psum)
  );
  basic_PE PE_Array_26_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_24_clock),
    .reset(PE_Array_26_24_reset),
    .io_in_activate(PE_Array_26_24_io_in_activate),
    .io_in_weight(PE_Array_26_24_io_in_weight),
    .io_in_psum(PE_Array_26_24_io_in_psum),
    .io_in_flow(PE_Array_26_24_io_in_flow),
    .io_in_shift(PE_Array_26_24_io_in_shift),
    .io_out_activate(PE_Array_26_24_io_out_activate),
    .io_out_weight(PE_Array_26_24_io_out_weight),
    .io_out_psum(PE_Array_26_24_io_out_psum)
  );
  basic_PE PE_Array_26_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_25_clock),
    .reset(PE_Array_26_25_reset),
    .io_in_activate(PE_Array_26_25_io_in_activate),
    .io_in_weight(PE_Array_26_25_io_in_weight),
    .io_in_psum(PE_Array_26_25_io_in_psum),
    .io_in_flow(PE_Array_26_25_io_in_flow),
    .io_in_shift(PE_Array_26_25_io_in_shift),
    .io_out_activate(PE_Array_26_25_io_out_activate),
    .io_out_weight(PE_Array_26_25_io_out_weight),
    .io_out_psum(PE_Array_26_25_io_out_psum)
  );
  basic_PE PE_Array_26_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_26_clock),
    .reset(PE_Array_26_26_reset),
    .io_in_activate(PE_Array_26_26_io_in_activate),
    .io_in_weight(PE_Array_26_26_io_in_weight),
    .io_in_psum(PE_Array_26_26_io_in_psum),
    .io_in_flow(PE_Array_26_26_io_in_flow),
    .io_in_shift(PE_Array_26_26_io_in_shift),
    .io_out_activate(PE_Array_26_26_io_out_activate),
    .io_out_weight(PE_Array_26_26_io_out_weight),
    .io_out_psum(PE_Array_26_26_io_out_psum)
  );
  basic_PE PE_Array_26_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_27_clock),
    .reset(PE_Array_26_27_reset),
    .io_in_activate(PE_Array_26_27_io_in_activate),
    .io_in_weight(PE_Array_26_27_io_in_weight),
    .io_in_psum(PE_Array_26_27_io_in_psum),
    .io_in_flow(PE_Array_26_27_io_in_flow),
    .io_in_shift(PE_Array_26_27_io_in_shift),
    .io_out_activate(PE_Array_26_27_io_out_activate),
    .io_out_weight(PE_Array_26_27_io_out_weight),
    .io_out_psum(PE_Array_26_27_io_out_psum)
  );
  basic_PE PE_Array_26_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_28_clock),
    .reset(PE_Array_26_28_reset),
    .io_in_activate(PE_Array_26_28_io_in_activate),
    .io_in_weight(PE_Array_26_28_io_in_weight),
    .io_in_psum(PE_Array_26_28_io_in_psum),
    .io_in_flow(PE_Array_26_28_io_in_flow),
    .io_in_shift(PE_Array_26_28_io_in_shift),
    .io_out_activate(PE_Array_26_28_io_out_activate),
    .io_out_weight(PE_Array_26_28_io_out_weight),
    .io_out_psum(PE_Array_26_28_io_out_psum)
  );
  basic_PE PE_Array_26_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_29_clock),
    .reset(PE_Array_26_29_reset),
    .io_in_activate(PE_Array_26_29_io_in_activate),
    .io_in_weight(PE_Array_26_29_io_in_weight),
    .io_in_psum(PE_Array_26_29_io_in_psum),
    .io_in_flow(PE_Array_26_29_io_in_flow),
    .io_in_shift(PE_Array_26_29_io_in_shift),
    .io_out_activate(PE_Array_26_29_io_out_activate),
    .io_out_weight(PE_Array_26_29_io_out_weight),
    .io_out_psum(PE_Array_26_29_io_out_psum)
  );
  basic_PE PE_Array_26_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_30_clock),
    .reset(PE_Array_26_30_reset),
    .io_in_activate(PE_Array_26_30_io_in_activate),
    .io_in_weight(PE_Array_26_30_io_in_weight),
    .io_in_psum(PE_Array_26_30_io_in_psum),
    .io_in_flow(PE_Array_26_30_io_in_flow),
    .io_in_shift(PE_Array_26_30_io_in_shift),
    .io_out_activate(PE_Array_26_30_io_out_activate),
    .io_out_weight(PE_Array_26_30_io_out_weight),
    .io_out_psum(PE_Array_26_30_io_out_psum)
  );
  basic_PE PE_Array_26_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_26_31_clock),
    .reset(PE_Array_26_31_reset),
    .io_in_activate(PE_Array_26_31_io_in_activate),
    .io_in_weight(PE_Array_26_31_io_in_weight),
    .io_in_psum(PE_Array_26_31_io_in_psum),
    .io_in_flow(PE_Array_26_31_io_in_flow),
    .io_in_shift(PE_Array_26_31_io_in_shift),
    .io_out_activate(PE_Array_26_31_io_out_activate),
    .io_out_weight(PE_Array_26_31_io_out_weight),
    .io_out_psum(PE_Array_26_31_io_out_psum)
  );
  basic_PE PE_Array_27_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_0_clock),
    .reset(PE_Array_27_0_reset),
    .io_in_activate(PE_Array_27_0_io_in_activate),
    .io_in_weight(PE_Array_27_0_io_in_weight),
    .io_in_psum(PE_Array_27_0_io_in_psum),
    .io_in_flow(PE_Array_27_0_io_in_flow),
    .io_in_shift(PE_Array_27_0_io_in_shift),
    .io_out_activate(PE_Array_27_0_io_out_activate),
    .io_out_weight(PE_Array_27_0_io_out_weight),
    .io_out_psum(PE_Array_27_0_io_out_psum)
  );
  basic_PE PE_Array_27_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_1_clock),
    .reset(PE_Array_27_1_reset),
    .io_in_activate(PE_Array_27_1_io_in_activate),
    .io_in_weight(PE_Array_27_1_io_in_weight),
    .io_in_psum(PE_Array_27_1_io_in_psum),
    .io_in_flow(PE_Array_27_1_io_in_flow),
    .io_in_shift(PE_Array_27_1_io_in_shift),
    .io_out_activate(PE_Array_27_1_io_out_activate),
    .io_out_weight(PE_Array_27_1_io_out_weight),
    .io_out_psum(PE_Array_27_1_io_out_psum)
  );
  basic_PE PE_Array_27_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_2_clock),
    .reset(PE_Array_27_2_reset),
    .io_in_activate(PE_Array_27_2_io_in_activate),
    .io_in_weight(PE_Array_27_2_io_in_weight),
    .io_in_psum(PE_Array_27_2_io_in_psum),
    .io_in_flow(PE_Array_27_2_io_in_flow),
    .io_in_shift(PE_Array_27_2_io_in_shift),
    .io_out_activate(PE_Array_27_2_io_out_activate),
    .io_out_weight(PE_Array_27_2_io_out_weight),
    .io_out_psum(PE_Array_27_2_io_out_psum)
  );
  basic_PE PE_Array_27_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_3_clock),
    .reset(PE_Array_27_3_reset),
    .io_in_activate(PE_Array_27_3_io_in_activate),
    .io_in_weight(PE_Array_27_3_io_in_weight),
    .io_in_psum(PE_Array_27_3_io_in_psum),
    .io_in_flow(PE_Array_27_3_io_in_flow),
    .io_in_shift(PE_Array_27_3_io_in_shift),
    .io_out_activate(PE_Array_27_3_io_out_activate),
    .io_out_weight(PE_Array_27_3_io_out_weight),
    .io_out_psum(PE_Array_27_3_io_out_psum)
  );
  basic_PE PE_Array_27_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_4_clock),
    .reset(PE_Array_27_4_reset),
    .io_in_activate(PE_Array_27_4_io_in_activate),
    .io_in_weight(PE_Array_27_4_io_in_weight),
    .io_in_psum(PE_Array_27_4_io_in_psum),
    .io_in_flow(PE_Array_27_4_io_in_flow),
    .io_in_shift(PE_Array_27_4_io_in_shift),
    .io_out_activate(PE_Array_27_4_io_out_activate),
    .io_out_weight(PE_Array_27_4_io_out_weight),
    .io_out_psum(PE_Array_27_4_io_out_psum)
  );
  basic_PE PE_Array_27_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_5_clock),
    .reset(PE_Array_27_5_reset),
    .io_in_activate(PE_Array_27_5_io_in_activate),
    .io_in_weight(PE_Array_27_5_io_in_weight),
    .io_in_psum(PE_Array_27_5_io_in_psum),
    .io_in_flow(PE_Array_27_5_io_in_flow),
    .io_in_shift(PE_Array_27_5_io_in_shift),
    .io_out_activate(PE_Array_27_5_io_out_activate),
    .io_out_weight(PE_Array_27_5_io_out_weight),
    .io_out_psum(PE_Array_27_5_io_out_psum)
  );
  basic_PE PE_Array_27_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_6_clock),
    .reset(PE_Array_27_6_reset),
    .io_in_activate(PE_Array_27_6_io_in_activate),
    .io_in_weight(PE_Array_27_6_io_in_weight),
    .io_in_psum(PE_Array_27_6_io_in_psum),
    .io_in_flow(PE_Array_27_6_io_in_flow),
    .io_in_shift(PE_Array_27_6_io_in_shift),
    .io_out_activate(PE_Array_27_6_io_out_activate),
    .io_out_weight(PE_Array_27_6_io_out_weight),
    .io_out_psum(PE_Array_27_6_io_out_psum)
  );
  basic_PE PE_Array_27_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_7_clock),
    .reset(PE_Array_27_7_reset),
    .io_in_activate(PE_Array_27_7_io_in_activate),
    .io_in_weight(PE_Array_27_7_io_in_weight),
    .io_in_psum(PE_Array_27_7_io_in_psum),
    .io_in_flow(PE_Array_27_7_io_in_flow),
    .io_in_shift(PE_Array_27_7_io_in_shift),
    .io_out_activate(PE_Array_27_7_io_out_activate),
    .io_out_weight(PE_Array_27_7_io_out_weight),
    .io_out_psum(PE_Array_27_7_io_out_psum)
  );
  basic_PE PE_Array_27_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_8_clock),
    .reset(PE_Array_27_8_reset),
    .io_in_activate(PE_Array_27_8_io_in_activate),
    .io_in_weight(PE_Array_27_8_io_in_weight),
    .io_in_psum(PE_Array_27_8_io_in_psum),
    .io_in_flow(PE_Array_27_8_io_in_flow),
    .io_in_shift(PE_Array_27_8_io_in_shift),
    .io_out_activate(PE_Array_27_8_io_out_activate),
    .io_out_weight(PE_Array_27_8_io_out_weight),
    .io_out_psum(PE_Array_27_8_io_out_psum)
  );
  basic_PE PE_Array_27_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_9_clock),
    .reset(PE_Array_27_9_reset),
    .io_in_activate(PE_Array_27_9_io_in_activate),
    .io_in_weight(PE_Array_27_9_io_in_weight),
    .io_in_psum(PE_Array_27_9_io_in_psum),
    .io_in_flow(PE_Array_27_9_io_in_flow),
    .io_in_shift(PE_Array_27_9_io_in_shift),
    .io_out_activate(PE_Array_27_9_io_out_activate),
    .io_out_weight(PE_Array_27_9_io_out_weight),
    .io_out_psum(PE_Array_27_9_io_out_psum)
  );
  basic_PE PE_Array_27_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_10_clock),
    .reset(PE_Array_27_10_reset),
    .io_in_activate(PE_Array_27_10_io_in_activate),
    .io_in_weight(PE_Array_27_10_io_in_weight),
    .io_in_psum(PE_Array_27_10_io_in_psum),
    .io_in_flow(PE_Array_27_10_io_in_flow),
    .io_in_shift(PE_Array_27_10_io_in_shift),
    .io_out_activate(PE_Array_27_10_io_out_activate),
    .io_out_weight(PE_Array_27_10_io_out_weight),
    .io_out_psum(PE_Array_27_10_io_out_psum)
  );
  basic_PE PE_Array_27_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_11_clock),
    .reset(PE_Array_27_11_reset),
    .io_in_activate(PE_Array_27_11_io_in_activate),
    .io_in_weight(PE_Array_27_11_io_in_weight),
    .io_in_psum(PE_Array_27_11_io_in_psum),
    .io_in_flow(PE_Array_27_11_io_in_flow),
    .io_in_shift(PE_Array_27_11_io_in_shift),
    .io_out_activate(PE_Array_27_11_io_out_activate),
    .io_out_weight(PE_Array_27_11_io_out_weight),
    .io_out_psum(PE_Array_27_11_io_out_psum)
  );
  basic_PE PE_Array_27_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_12_clock),
    .reset(PE_Array_27_12_reset),
    .io_in_activate(PE_Array_27_12_io_in_activate),
    .io_in_weight(PE_Array_27_12_io_in_weight),
    .io_in_psum(PE_Array_27_12_io_in_psum),
    .io_in_flow(PE_Array_27_12_io_in_flow),
    .io_in_shift(PE_Array_27_12_io_in_shift),
    .io_out_activate(PE_Array_27_12_io_out_activate),
    .io_out_weight(PE_Array_27_12_io_out_weight),
    .io_out_psum(PE_Array_27_12_io_out_psum)
  );
  basic_PE PE_Array_27_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_13_clock),
    .reset(PE_Array_27_13_reset),
    .io_in_activate(PE_Array_27_13_io_in_activate),
    .io_in_weight(PE_Array_27_13_io_in_weight),
    .io_in_psum(PE_Array_27_13_io_in_psum),
    .io_in_flow(PE_Array_27_13_io_in_flow),
    .io_in_shift(PE_Array_27_13_io_in_shift),
    .io_out_activate(PE_Array_27_13_io_out_activate),
    .io_out_weight(PE_Array_27_13_io_out_weight),
    .io_out_psum(PE_Array_27_13_io_out_psum)
  );
  basic_PE PE_Array_27_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_14_clock),
    .reset(PE_Array_27_14_reset),
    .io_in_activate(PE_Array_27_14_io_in_activate),
    .io_in_weight(PE_Array_27_14_io_in_weight),
    .io_in_psum(PE_Array_27_14_io_in_psum),
    .io_in_flow(PE_Array_27_14_io_in_flow),
    .io_in_shift(PE_Array_27_14_io_in_shift),
    .io_out_activate(PE_Array_27_14_io_out_activate),
    .io_out_weight(PE_Array_27_14_io_out_weight),
    .io_out_psum(PE_Array_27_14_io_out_psum)
  );
  basic_PE PE_Array_27_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_15_clock),
    .reset(PE_Array_27_15_reset),
    .io_in_activate(PE_Array_27_15_io_in_activate),
    .io_in_weight(PE_Array_27_15_io_in_weight),
    .io_in_psum(PE_Array_27_15_io_in_psum),
    .io_in_flow(PE_Array_27_15_io_in_flow),
    .io_in_shift(PE_Array_27_15_io_in_shift),
    .io_out_activate(PE_Array_27_15_io_out_activate),
    .io_out_weight(PE_Array_27_15_io_out_weight),
    .io_out_psum(PE_Array_27_15_io_out_psum)
  );
  basic_PE PE_Array_27_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_16_clock),
    .reset(PE_Array_27_16_reset),
    .io_in_activate(PE_Array_27_16_io_in_activate),
    .io_in_weight(PE_Array_27_16_io_in_weight),
    .io_in_psum(PE_Array_27_16_io_in_psum),
    .io_in_flow(PE_Array_27_16_io_in_flow),
    .io_in_shift(PE_Array_27_16_io_in_shift),
    .io_out_activate(PE_Array_27_16_io_out_activate),
    .io_out_weight(PE_Array_27_16_io_out_weight),
    .io_out_psum(PE_Array_27_16_io_out_psum)
  );
  basic_PE PE_Array_27_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_17_clock),
    .reset(PE_Array_27_17_reset),
    .io_in_activate(PE_Array_27_17_io_in_activate),
    .io_in_weight(PE_Array_27_17_io_in_weight),
    .io_in_psum(PE_Array_27_17_io_in_psum),
    .io_in_flow(PE_Array_27_17_io_in_flow),
    .io_in_shift(PE_Array_27_17_io_in_shift),
    .io_out_activate(PE_Array_27_17_io_out_activate),
    .io_out_weight(PE_Array_27_17_io_out_weight),
    .io_out_psum(PE_Array_27_17_io_out_psum)
  );
  basic_PE PE_Array_27_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_18_clock),
    .reset(PE_Array_27_18_reset),
    .io_in_activate(PE_Array_27_18_io_in_activate),
    .io_in_weight(PE_Array_27_18_io_in_weight),
    .io_in_psum(PE_Array_27_18_io_in_psum),
    .io_in_flow(PE_Array_27_18_io_in_flow),
    .io_in_shift(PE_Array_27_18_io_in_shift),
    .io_out_activate(PE_Array_27_18_io_out_activate),
    .io_out_weight(PE_Array_27_18_io_out_weight),
    .io_out_psum(PE_Array_27_18_io_out_psum)
  );
  basic_PE PE_Array_27_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_19_clock),
    .reset(PE_Array_27_19_reset),
    .io_in_activate(PE_Array_27_19_io_in_activate),
    .io_in_weight(PE_Array_27_19_io_in_weight),
    .io_in_psum(PE_Array_27_19_io_in_psum),
    .io_in_flow(PE_Array_27_19_io_in_flow),
    .io_in_shift(PE_Array_27_19_io_in_shift),
    .io_out_activate(PE_Array_27_19_io_out_activate),
    .io_out_weight(PE_Array_27_19_io_out_weight),
    .io_out_psum(PE_Array_27_19_io_out_psum)
  );
  basic_PE PE_Array_27_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_20_clock),
    .reset(PE_Array_27_20_reset),
    .io_in_activate(PE_Array_27_20_io_in_activate),
    .io_in_weight(PE_Array_27_20_io_in_weight),
    .io_in_psum(PE_Array_27_20_io_in_psum),
    .io_in_flow(PE_Array_27_20_io_in_flow),
    .io_in_shift(PE_Array_27_20_io_in_shift),
    .io_out_activate(PE_Array_27_20_io_out_activate),
    .io_out_weight(PE_Array_27_20_io_out_weight),
    .io_out_psum(PE_Array_27_20_io_out_psum)
  );
  basic_PE PE_Array_27_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_21_clock),
    .reset(PE_Array_27_21_reset),
    .io_in_activate(PE_Array_27_21_io_in_activate),
    .io_in_weight(PE_Array_27_21_io_in_weight),
    .io_in_psum(PE_Array_27_21_io_in_psum),
    .io_in_flow(PE_Array_27_21_io_in_flow),
    .io_in_shift(PE_Array_27_21_io_in_shift),
    .io_out_activate(PE_Array_27_21_io_out_activate),
    .io_out_weight(PE_Array_27_21_io_out_weight),
    .io_out_psum(PE_Array_27_21_io_out_psum)
  );
  basic_PE PE_Array_27_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_22_clock),
    .reset(PE_Array_27_22_reset),
    .io_in_activate(PE_Array_27_22_io_in_activate),
    .io_in_weight(PE_Array_27_22_io_in_weight),
    .io_in_psum(PE_Array_27_22_io_in_psum),
    .io_in_flow(PE_Array_27_22_io_in_flow),
    .io_in_shift(PE_Array_27_22_io_in_shift),
    .io_out_activate(PE_Array_27_22_io_out_activate),
    .io_out_weight(PE_Array_27_22_io_out_weight),
    .io_out_psum(PE_Array_27_22_io_out_psum)
  );
  basic_PE PE_Array_27_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_23_clock),
    .reset(PE_Array_27_23_reset),
    .io_in_activate(PE_Array_27_23_io_in_activate),
    .io_in_weight(PE_Array_27_23_io_in_weight),
    .io_in_psum(PE_Array_27_23_io_in_psum),
    .io_in_flow(PE_Array_27_23_io_in_flow),
    .io_in_shift(PE_Array_27_23_io_in_shift),
    .io_out_activate(PE_Array_27_23_io_out_activate),
    .io_out_weight(PE_Array_27_23_io_out_weight),
    .io_out_psum(PE_Array_27_23_io_out_psum)
  );
  basic_PE PE_Array_27_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_24_clock),
    .reset(PE_Array_27_24_reset),
    .io_in_activate(PE_Array_27_24_io_in_activate),
    .io_in_weight(PE_Array_27_24_io_in_weight),
    .io_in_psum(PE_Array_27_24_io_in_psum),
    .io_in_flow(PE_Array_27_24_io_in_flow),
    .io_in_shift(PE_Array_27_24_io_in_shift),
    .io_out_activate(PE_Array_27_24_io_out_activate),
    .io_out_weight(PE_Array_27_24_io_out_weight),
    .io_out_psum(PE_Array_27_24_io_out_psum)
  );
  basic_PE PE_Array_27_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_25_clock),
    .reset(PE_Array_27_25_reset),
    .io_in_activate(PE_Array_27_25_io_in_activate),
    .io_in_weight(PE_Array_27_25_io_in_weight),
    .io_in_psum(PE_Array_27_25_io_in_psum),
    .io_in_flow(PE_Array_27_25_io_in_flow),
    .io_in_shift(PE_Array_27_25_io_in_shift),
    .io_out_activate(PE_Array_27_25_io_out_activate),
    .io_out_weight(PE_Array_27_25_io_out_weight),
    .io_out_psum(PE_Array_27_25_io_out_psum)
  );
  basic_PE PE_Array_27_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_26_clock),
    .reset(PE_Array_27_26_reset),
    .io_in_activate(PE_Array_27_26_io_in_activate),
    .io_in_weight(PE_Array_27_26_io_in_weight),
    .io_in_psum(PE_Array_27_26_io_in_psum),
    .io_in_flow(PE_Array_27_26_io_in_flow),
    .io_in_shift(PE_Array_27_26_io_in_shift),
    .io_out_activate(PE_Array_27_26_io_out_activate),
    .io_out_weight(PE_Array_27_26_io_out_weight),
    .io_out_psum(PE_Array_27_26_io_out_psum)
  );
  basic_PE PE_Array_27_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_27_clock),
    .reset(PE_Array_27_27_reset),
    .io_in_activate(PE_Array_27_27_io_in_activate),
    .io_in_weight(PE_Array_27_27_io_in_weight),
    .io_in_psum(PE_Array_27_27_io_in_psum),
    .io_in_flow(PE_Array_27_27_io_in_flow),
    .io_in_shift(PE_Array_27_27_io_in_shift),
    .io_out_activate(PE_Array_27_27_io_out_activate),
    .io_out_weight(PE_Array_27_27_io_out_weight),
    .io_out_psum(PE_Array_27_27_io_out_psum)
  );
  basic_PE PE_Array_27_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_28_clock),
    .reset(PE_Array_27_28_reset),
    .io_in_activate(PE_Array_27_28_io_in_activate),
    .io_in_weight(PE_Array_27_28_io_in_weight),
    .io_in_psum(PE_Array_27_28_io_in_psum),
    .io_in_flow(PE_Array_27_28_io_in_flow),
    .io_in_shift(PE_Array_27_28_io_in_shift),
    .io_out_activate(PE_Array_27_28_io_out_activate),
    .io_out_weight(PE_Array_27_28_io_out_weight),
    .io_out_psum(PE_Array_27_28_io_out_psum)
  );
  basic_PE PE_Array_27_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_29_clock),
    .reset(PE_Array_27_29_reset),
    .io_in_activate(PE_Array_27_29_io_in_activate),
    .io_in_weight(PE_Array_27_29_io_in_weight),
    .io_in_psum(PE_Array_27_29_io_in_psum),
    .io_in_flow(PE_Array_27_29_io_in_flow),
    .io_in_shift(PE_Array_27_29_io_in_shift),
    .io_out_activate(PE_Array_27_29_io_out_activate),
    .io_out_weight(PE_Array_27_29_io_out_weight),
    .io_out_psum(PE_Array_27_29_io_out_psum)
  );
  basic_PE PE_Array_27_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_30_clock),
    .reset(PE_Array_27_30_reset),
    .io_in_activate(PE_Array_27_30_io_in_activate),
    .io_in_weight(PE_Array_27_30_io_in_weight),
    .io_in_psum(PE_Array_27_30_io_in_psum),
    .io_in_flow(PE_Array_27_30_io_in_flow),
    .io_in_shift(PE_Array_27_30_io_in_shift),
    .io_out_activate(PE_Array_27_30_io_out_activate),
    .io_out_weight(PE_Array_27_30_io_out_weight),
    .io_out_psum(PE_Array_27_30_io_out_psum)
  );
  basic_PE PE_Array_27_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_27_31_clock),
    .reset(PE_Array_27_31_reset),
    .io_in_activate(PE_Array_27_31_io_in_activate),
    .io_in_weight(PE_Array_27_31_io_in_weight),
    .io_in_psum(PE_Array_27_31_io_in_psum),
    .io_in_flow(PE_Array_27_31_io_in_flow),
    .io_in_shift(PE_Array_27_31_io_in_shift),
    .io_out_activate(PE_Array_27_31_io_out_activate),
    .io_out_weight(PE_Array_27_31_io_out_weight),
    .io_out_psum(PE_Array_27_31_io_out_psum)
  );
  basic_PE PE_Array_28_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_0_clock),
    .reset(PE_Array_28_0_reset),
    .io_in_activate(PE_Array_28_0_io_in_activate),
    .io_in_weight(PE_Array_28_0_io_in_weight),
    .io_in_psum(PE_Array_28_0_io_in_psum),
    .io_in_flow(PE_Array_28_0_io_in_flow),
    .io_in_shift(PE_Array_28_0_io_in_shift),
    .io_out_activate(PE_Array_28_0_io_out_activate),
    .io_out_weight(PE_Array_28_0_io_out_weight),
    .io_out_psum(PE_Array_28_0_io_out_psum)
  );
  basic_PE PE_Array_28_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_1_clock),
    .reset(PE_Array_28_1_reset),
    .io_in_activate(PE_Array_28_1_io_in_activate),
    .io_in_weight(PE_Array_28_1_io_in_weight),
    .io_in_psum(PE_Array_28_1_io_in_psum),
    .io_in_flow(PE_Array_28_1_io_in_flow),
    .io_in_shift(PE_Array_28_1_io_in_shift),
    .io_out_activate(PE_Array_28_1_io_out_activate),
    .io_out_weight(PE_Array_28_1_io_out_weight),
    .io_out_psum(PE_Array_28_1_io_out_psum)
  );
  basic_PE PE_Array_28_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_2_clock),
    .reset(PE_Array_28_2_reset),
    .io_in_activate(PE_Array_28_2_io_in_activate),
    .io_in_weight(PE_Array_28_2_io_in_weight),
    .io_in_psum(PE_Array_28_2_io_in_psum),
    .io_in_flow(PE_Array_28_2_io_in_flow),
    .io_in_shift(PE_Array_28_2_io_in_shift),
    .io_out_activate(PE_Array_28_2_io_out_activate),
    .io_out_weight(PE_Array_28_2_io_out_weight),
    .io_out_psum(PE_Array_28_2_io_out_psum)
  );
  basic_PE PE_Array_28_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_3_clock),
    .reset(PE_Array_28_3_reset),
    .io_in_activate(PE_Array_28_3_io_in_activate),
    .io_in_weight(PE_Array_28_3_io_in_weight),
    .io_in_psum(PE_Array_28_3_io_in_psum),
    .io_in_flow(PE_Array_28_3_io_in_flow),
    .io_in_shift(PE_Array_28_3_io_in_shift),
    .io_out_activate(PE_Array_28_3_io_out_activate),
    .io_out_weight(PE_Array_28_3_io_out_weight),
    .io_out_psum(PE_Array_28_3_io_out_psum)
  );
  basic_PE PE_Array_28_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_4_clock),
    .reset(PE_Array_28_4_reset),
    .io_in_activate(PE_Array_28_4_io_in_activate),
    .io_in_weight(PE_Array_28_4_io_in_weight),
    .io_in_psum(PE_Array_28_4_io_in_psum),
    .io_in_flow(PE_Array_28_4_io_in_flow),
    .io_in_shift(PE_Array_28_4_io_in_shift),
    .io_out_activate(PE_Array_28_4_io_out_activate),
    .io_out_weight(PE_Array_28_4_io_out_weight),
    .io_out_psum(PE_Array_28_4_io_out_psum)
  );
  basic_PE PE_Array_28_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_5_clock),
    .reset(PE_Array_28_5_reset),
    .io_in_activate(PE_Array_28_5_io_in_activate),
    .io_in_weight(PE_Array_28_5_io_in_weight),
    .io_in_psum(PE_Array_28_5_io_in_psum),
    .io_in_flow(PE_Array_28_5_io_in_flow),
    .io_in_shift(PE_Array_28_5_io_in_shift),
    .io_out_activate(PE_Array_28_5_io_out_activate),
    .io_out_weight(PE_Array_28_5_io_out_weight),
    .io_out_psum(PE_Array_28_5_io_out_psum)
  );
  basic_PE PE_Array_28_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_6_clock),
    .reset(PE_Array_28_6_reset),
    .io_in_activate(PE_Array_28_6_io_in_activate),
    .io_in_weight(PE_Array_28_6_io_in_weight),
    .io_in_psum(PE_Array_28_6_io_in_psum),
    .io_in_flow(PE_Array_28_6_io_in_flow),
    .io_in_shift(PE_Array_28_6_io_in_shift),
    .io_out_activate(PE_Array_28_6_io_out_activate),
    .io_out_weight(PE_Array_28_6_io_out_weight),
    .io_out_psum(PE_Array_28_6_io_out_psum)
  );
  basic_PE PE_Array_28_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_7_clock),
    .reset(PE_Array_28_7_reset),
    .io_in_activate(PE_Array_28_7_io_in_activate),
    .io_in_weight(PE_Array_28_7_io_in_weight),
    .io_in_psum(PE_Array_28_7_io_in_psum),
    .io_in_flow(PE_Array_28_7_io_in_flow),
    .io_in_shift(PE_Array_28_7_io_in_shift),
    .io_out_activate(PE_Array_28_7_io_out_activate),
    .io_out_weight(PE_Array_28_7_io_out_weight),
    .io_out_psum(PE_Array_28_7_io_out_psum)
  );
  basic_PE PE_Array_28_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_8_clock),
    .reset(PE_Array_28_8_reset),
    .io_in_activate(PE_Array_28_8_io_in_activate),
    .io_in_weight(PE_Array_28_8_io_in_weight),
    .io_in_psum(PE_Array_28_8_io_in_psum),
    .io_in_flow(PE_Array_28_8_io_in_flow),
    .io_in_shift(PE_Array_28_8_io_in_shift),
    .io_out_activate(PE_Array_28_8_io_out_activate),
    .io_out_weight(PE_Array_28_8_io_out_weight),
    .io_out_psum(PE_Array_28_8_io_out_psum)
  );
  basic_PE PE_Array_28_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_9_clock),
    .reset(PE_Array_28_9_reset),
    .io_in_activate(PE_Array_28_9_io_in_activate),
    .io_in_weight(PE_Array_28_9_io_in_weight),
    .io_in_psum(PE_Array_28_9_io_in_psum),
    .io_in_flow(PE_Array_28_9_io_in_flow),
    .io_in_shift(PE_Array_28_9_io_in_shift),
    .io_out_activate(PE_Array_28_9_io_out_activate),
    .io_out_weight(PE_Array_28_9_io_out_weight),
    .io_out_psum(PE_Array_28_9_io_out_psum)
  );
  basic_PE PE_Array_28_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_10_clock),
    .reset(PE_Array_28_10_reset),
    .io_in_activate(PE_Array_28_10_io_in_activate),
    .io_in_weight(PE_Array_28_10_io_in_weight),
    .io_in_psum(PE_Array_28_10_io_in_psum),
    .io_in_flow(PE_Array_28_10_io_in_flow),
    .io_in_shift(PE_Array_28_10_io_in_shift),
    .io_out_activate(PE_Array_28_10_io_out_activate),
    .io_out_weight(PE_Array_28_10_io_out_weight),
    .io_out_psum(PE_Array_28_10_io_out_psum)
  );
  basic_PE PE_Array_28_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_11_clock),
    .reset(PE_Array_28_11_reset),
    .io_in_activate(PE_Array_28_11_io_in_activate),
    .io_in_weight(PE_Array_28_11_io_in_weight),
    .io_in_psum(PE_Array_28_11_io_in_psum),
    .io_in_flow(PE_Array_28_11_io_in_flow),
    .io_in_shift(PE_Array_28_11_io_in_shift),
    .io_out_activate(PE_Array_28_11_io_out_activate),
    .io_out_weight(PE_Array_28_11_io_out_weight),
    .io_out_psum(PE_Array_28_11_io_out_psum)
  );
  basic_PE PE_Array_28_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_12_clock),
    .reset(PE_Array_28_12_reset),
    .io_in_activate(PE_Array_28_12_io_in_activate),
    .io_in_weight(PE_Array_28_12_io_in_weight),
    .io_in_psum(PE_Array_28_12_io_in_psum),
    .io_in_flow(PE_Array_28_12_io_in_flow),
    .io_in_shift(PE_Array_28_12_io_in_shift),
    .io_out_activate(PE_Array_28_12_io_out_activate),
    .io_out_weight(PE_Array_28_12_io_out_weight),
    .io_out_psum(PE_Array_28_12_io_out_psum)
  );
  basic_PE PE_Array_28_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_13_clock),
    .reset(PE_Array_28_13_reset),
    .io_in_activate(PE_Array_28_13_io_in_activate),
    .io_in_weight(PE_Array_28_13_io_in_weight),
    .io_in_psum(PE_Array_28_13_io_in_psum),
    .io_in_flow(PE_Array_28_13_io_in_flow),
    .io_in_shift(PE_Array_28_13_io_in_shift),
    .io_out_activate(PE_Array_28_13_io_out_activate),
    .io_out_weight(PE_Array_28_13_io_out_weight),
    .io_out_psum(PE_Array_28_13_io_out_psum)
  );
  basic_PE PE_Array_28_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_14_clock),
    .reset(PE_Array_28_14_reset),
    .io_in_activate(PE_Array_28_14_io_in_activate),
    .io_in_weight(PE_Array_28_14_io_in_weight),
    .io_in_psum(PE_Array_28_14_io_in_psum),
    .io_in_flow(PE_Array_28_14_io_in_flow),
    .io_in_shift(PE_Array_28_14_io_in_shift),
    .io_out_activate(PE_Array_28_14_io_out_activate),
    .io_out_weight(PE_Array_28_14_io_out_weight),
    .io_out_psum(PE_Array_28_14_io_out_psum)
  );
  basic_PE PE_Array_28_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_15_clock),
    .reset(PE_Array_28_15_reset),
    .io_in_activate(PE_Array_28_15_io_in_activate),
    .io_in_weight(PE_Array_28_15_io_in_weight),
    .io_in_psum(PE_Array_28_15_io_in_psum),
    .io_in_flow(PE_Array_28_15_io_in_flow),
    .io_in_shift(PE_Array_28_15_io_in_shift),
    .io_out_activate(PE_Array_28_15_io_out_activate),
    .io_out_weight(PE_Array_28_15_io_out_weight),
    .io_out_psum(PE_Array_28_15_io_out_psum)
  );
  basic_PE PE_Array_28_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_16_clock),
    .reset(PE_Array_28_16_reset),
    .io_in_activate(PE_Array_28_16_io_in_activate),
    .io_in_weight(PE_Array_28_16_io_in_weight),
    .io_in_psum(PE_Array_28_16_io_in_psum),
    .io_in_flow(PE_Array_28_16_io_in_flow),
    .io_in_shift(PE_Array_28_16_io_in_shift),
    .io_out_activate(PE_Array_28_16_io_out_activate),
    .io_out_weight(PE_Array_28_16_io_out_weight),
    .io_out_psum(PE_Array_28_16_io_out_psum)
  );
  basic_PE PE_Array_28_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_17_clock),
    .reset(PE_Array_28_17_reset),
    .io_in_activate(PE_Array_28_17_io_in_activate),
    .io_in_weight(PE_Array_28_17_io_in_weight),
    .io_in_psum(PE_Array_28_17_io_in_psum),
    .io_in_flow(PE_Array_28_17_io_in_flow),
    .io_in_shift(PE_Array_28_17_io_in_shift),
    .io_out_activate(PE_Array_28_17_io_out_activate),
    .io_out_weight(PE_Array_28_17_io_out_weight),
    .io_out_psum(PE_Array_28_17_io_out_psum)
  );
  basic_PE PE_Array_28_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_18_clock),
    .reset(PE_Array_28_18_reset),
    .io_in_activate(PE_Array_28_18_io_in_activate),
    .io_in_weight(PE_Array_28_18_io_in_weight),
    .io_in_psum(PE_Array_28_18_io_in_psum),
    .io_in_flow(PE_Array_28_18_io_in_flow),
    .io_in_shift(PE_Array_28_18_io_in_shift),
    .io_out_activate(PE_Array_28_18_io_out_activate),
    .io_out_weight(PE_Array_28_18_io_out_weight),
    .io_out_psum(PE_Array_28_18_io_out_psum)
  );
  basic_PE PE_Array_28_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_19_clock),
    .reset(PE_Array_28_19_reset),
    .io_in_activate(PE_Array_28_19_io_in_activate),
    .io_in_weight(PE_Array_28_19_io_in_weight),
    .io_in_psum(PE_Array_28_19_io_in_psum),
    .io_in_flow(PE_Array_28_19_io_in_flow),
    .io_in_shift(PE_Array_28_19_io_in_shift),
    .io_out_activate(PE_Array_28_19_io_out_activate),
    .io_out_weight(PE_Array_28_19_io_out_weight),
    .io_out_psum(PE_Array_28_19_io_out_psum)
  );
  basic_PE PE_Array_28_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_20_clock),
    .reset(PE_Array_28_20_reset),
    .io_in_activate(PE_Array_28_20_io_in_activate),
    .io_in_weight(PE_Array_28_20_io_in_weight),
    .io_in_psum(PE_Array_28_20_io_in_psum),
    .io_in_flow(PE_Array_28_20_io_in_flow),
    .io_in_shift(PE_Array_28_20_io_in_shift),
    .io_out_activate(PE_Array_28_20_io_out_activate),
    .io_out_weight(PE_Array_28_20_io_out_weight),
    .io_out_psum(PE_Array_28_20_io_out_psum)
  );
  basic_PE PE_Array_28_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_21_clock),
    .reset(PE_Array_28_21_reset),
    .io_in_activate(PE_Array_28_21_io_in_activate),
    .io_in_weight(PE_Array_28_21_io_in_weight),
    .io_in_psum(PE_Array_28_21_io_in_psum),
    .io_in_flow(PE_Array_28_21_io_in_flow),
    .io_in_shift(PE_Array_28_21_io_in_shift),
    .io_out_activate(PE_Array_28_21_io_out_activate),
    .io_out_weight(PE_Array_28_21_io_out_weight),
    .io_out_psum(PE_Array_28_21_io_out_psum)
  );
  basic_PE PE_Array_28_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_22_clock),
    .reset(PE_Array_28_22_reset),
    .io_in_activate(PE_Array_28_22_io_in_activate),
    .io_in_weight(PE_Array_28_22_io_in_weight),
    .io_in_psum(PE_Array_28_22_io_in_psum),
    .io_in_flow(PE_Array_28_22_io_in_flow),
    .io_in_shift(PE_Array_28_22_io_in_shift),
    .io_out_activate(PE_Array_28_22_io_out_activate),
    .io_out_weight(PE_Array_28_22_io_out_weight),
    .io_out_psum(PE_Array_28_22_io_out_psum)
  );
  basic_PE PE_Array_28_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_23_clock),
    .reset(PE_Array_28_23_reset),
    .io_in_activate(PE_Array_28_23_io_in_activate),
    .io_in_weight(PE_Array_28_23_io_in_weight),
    .io_in_psum(PE_Array_28_23_io_in_psum),
    .io_in_flow(PE_Array_28_23_io_in_flow),
    .io_in_shift(PE_Array_28_23_io_in_shift),
    .io_out_activate(PE_Array_28_23_io_out_activate),
    .io_out_weight(PE_Array_28_23_io_out_weight),
    .io_out_psum(PE_Array_28_23_io_out_psum)
  );
  basic_PE PE_Array_28_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_24_clock),
    .reset(PE_Array_28_24_reset),
    .io_in_activate(PE_Array_28_24_io_in_activate),
    .io_in_weight(PE_Array_28_24_io_in_weight),
    .io_in_psum(PE_Array_28_24_io_in_psum),
    .io_in_flow(PE_Array_28_24_io_in_flow),
    .io_in_shift(PE_Array_28_24_io_in_shift),
    .io_out_activate(PE_Array_28_24_io_out_activate),
    .io_out_weight(PE_Array_28_24_io_out_weight),
    .io_out_psum(PE_Array_28_24_io_out_psum)
  );
  basic_PE PE_Array_28_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_25_clock),
    .reset(PE_Array_28_25_reset),
    .io_in_activate(PE_Array_28_25_io_in_activate),
    .io_in_weight(PE_Array_28_25_io_in_weight),
    .io_in_psum(PE_Array_28_25_io_in_psum),
    .io_in_flow(PE_Array_28_25_io_in_flow),
    .io_in_shift(PE_Array_28_25_io_in_shift),
    .io_out_activate(PE_Array_28_25_io_out_activate),
    .io_out_weight(PE_Array_28_25_io_out_weight),
    .io_out_psum(PE_Array_28_25_io_out_psum)
  );
  basic_PE PE_Array_28_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_26_clock),
    .reset(PE_Array_28_26_reset),
    .io_in_activate(PE_Array_28_26_io_in_activate),
    .io_in_weight(PE_Array_28_26_io_in_weight),
    .io_in_psum(PE_Array_28_26_io_in_psum),
    .io_in_flow(PE_Array_28_26_io_in_flow),
    .io_in_shift(PE_Array_28_26_io_in_shift),
    .io_out_activate(PE_Array_28_26_io_out_activate),
    .io_out_weight(PE_Array_28_26_io_out_weight),
    .io_out_psum(PE_Array_28_26_io_out_psum)
  );
  basic_PE PE_Array_28_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_27_clock),
    .reset(PE_Array_28_27_reset),
    .io_in_activate(PE_Array_28_27_io_in_activate),
    .io_in_weight(PE_Array_28_27_io_in_weight),
    .io_in_psum(PE_Array_28_27_io_in_psum),
    .io_in_flow(PE_Array_28_27_io_in_flow),
    .io_in_shift(PE_Array_28_27_io_in_shift),
    .io_out_activate(PE_Array_28_27_io_out_activate),
    .io_out_weight(PE_Array_28_27_io_out_weight),
    .io_out_psum(PE_Array_28_27_io_out_psum)
  );
  basic_PE PE_Array_28_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_28_clock),
    .reset(PE_Array_28_28_reset),
    .io_in_activate(PE_Array_28_28_io_in_activate),
    .io_in_weight(PE_Array_28_28_io_in_weight),
    .io_in_psum(PE_Array_28_28_io_in_psum),
    .io_in_flow(PE_Array_28_28_io_in_flow),
    .io_in_shift(PE_Array_28_28_io_in_shift),
    .io_out_activate(PE_Array_28_28_io_out_activate),
    .io_out_weight(PE_Array_28_28_io_out_weight),
    .io_out_psum(PE_Array_28_28_io_out_psum)
  );
  basic_PE PE_Array_28_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_29_clock),
    .reset(PE_Array_28_29_reset),
    .io_in_activate(PE_Array_28_29_io_in_activate),
    .io_in_weight(PE_Array_28_29_io_in_weight),
    .io_in_psum(PE_Array_28_29_io_in_psum),
    .io_in_flow(PE_Array_28_29_io_in_flow),
    .io_in_shift(PE_Array_28_29_io_in_shift),
    .io_out_activate(PE_Array_28_29_io_out_activate),
    .io_out_weight(PE_Array_28_29_io_out_weight),
    .io_out_psum(PE_Array_28_29_io_out_psum)
  );
  basic_PE PE_Array_28_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_30_clock),
    .reset(PE_Array_28_30_reset),
    .io_in_activate(PE_Array_28_30_io_in_activate),
    .io_in_weight(PE_Array_28_30_io_in_weight),
    .io_in_psum(PE_Array_28_30_io_in_psum),
    .io_in_flow(PE_Array_28_30_io_in_flow),
    .io_in_shift(PE_Array_28_30_io_in_shift),
    .io_out_activate(PE_Array_28_30_io_out_activate),
    .io_out_weight(PE_Array_28_30_io_out_weight),
    .io_out_psum(PE_Array_28_30_io_out_psum)
  );
  basic_PE PE_Array_28_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_28_31_clock),
    .reset(PE_Array_28_31_reset),
    .io_in_activate(PE_Array_28_31_io_in_activate),
    .io_in_weight(PE_Array_28_31_io_in_weight),
    .io_in_psum(PE_Array_28_31_io_in_psum),
    .io_in_flow(PE_Array_28_31_io_in_flow),
    .io_in_shift(PE_Array_28_31_io_in_shift),
    .io_out_activate(PE_Array_28_31_io_out_activate),
    .io_out_weight(PE_Array_28_31_io_out_weight),
    .io_out_psum(PE_Array_28_31_io_out_psum)
  );
  basic_PE PE_Array_29_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_0_clock),
    .reset(PE_Array_29_0_reset),
    .io_in_activate(PE_Array_29_0_io_in_activate),
    .io_in_weight(PE_Array_29_0_io_in_weight),
    .io_in_psum(PE_Array_29_0_io_in_psum),
    .io_in_flow(PE_Array_29_0_io_in_flow),
    .io_in_shift(PE_Array_29_0_io_in_shift),
    .io_out_activate(PE_Array_29_0_io_out_activate),
    .io_out_weight(PE_Array_29_0_io_out_weight),
    .io_out_psum(PE_Array_29_0_io_out_psum)
  );
  basic_PE PE_Array_29_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_1_clock),
    .reset(PE_Array_29_1_reset),
    .io_in_activate(PE_Array_29_1_io_in_activate),
    .io_in_weight(PE_Array_29_1_io_in_weight),
    .io_in_psum(PE_Array_29_1_io_in_psum),
    .io_in_flow(PE_Array_29_1_io_in_flow),
    .io_in_shift(PE_Array_29_1_io_in_shift),
    .io_out_activate(PE_Array_29_1_io_out_activate),
    .io_out_weight(PE_Array_29_1_io_out_weight),
    .io_out_psum(PE_Array_29_1_io_out_psum)
  );
  basic_PE PE_Array_29_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_2_clock),
    .reset(PE_Array_29_2_reset),
    .io_in_activate(PE_Array_29_2_io_in_activate),
    .io_in_weight(PE_Array_29_2_io_in_weight),
    .io_in_psum(PE_Array_29_2_io_in_psum),
    .io_in_flow(PE_Array_29_2_io_in_flow),
    .io_in_shift(PE_Array_29_2_io_in_shift),
    .io_out_activate(PE_Array_29_2_io_out_activate),
    .io_out_weight(PE_Array_29_2_io_out_weight),
    .io_out_psum(PE_Array_29_2_io_out_psum)
  );
  basic_PE PE_Array_29_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_3_clock),
    .reset(PE_Array_29_3_reset),
    .io_in_activate(PE_Array_29_3_io_in_activate),
    .io_in_weight(PE_Array_29_3_io_in_weight),
    .io_in_psum(PE_Array_29_3_io_in_psum),
    .io_in_flow(PE_Array_29_3_io_in_flow),
    .io_in_shift(PE_Array_29_3_io_in_shift),
    .io_out_activate(PE_Array_29_3_io_out_activate),
    .io_out_weight(PE_Array_29_3_io_out_weight),
    .io_out_psum(PE_Array_29_3_io_out_psum)
  );
  basic_PE PE_Array_29_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_4_clock),
    .reset(PE_Array_29_4_reset),
    .io_in_activate(PE_Array_29_4_io_in_activate),
    .io_in_weight(PE_Array_29_4_io_in_weight),
    .io_in_psum(PE_Array_29_4_io_in_psum),
    .io_in_flow(PE_Array_29_4_io_in_flow),
    .io_in_shift(PE_Array_29_4_io_in_shift),
    .io_out_activate(PE_Array_29_4_io_out_activate),
    .io_out_weight(PE_Array_29_4_io_out_weight),
    .io_out_psum(PE_Array_29_4_io_out_psum)
  );
  basic_PE PE_Array_29_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_5_clock),
    .reset(PE_Array_29_5_reset),
    .io_in_activate(PE_Array_29_5_io_in_activate),
    .io_in_weight(PE_Array_29_5_io_in_weight),
    .io_in_psum(PE_Array_29_5_io_in_psum),
    .io_in_flow(PE_Array_29_5_io_in_flow),
    .io_in_shift(PE_Array_29_5_io_in_shift),
    .io_out_activate(PE_Array_29_5_io_out_activate),
    .io_out_weight(PE_Array_29_5_io_out_weight),
    .io_out_psum(PE_Array_29_5_io_out_psum)
  );
  basic_PE PE_Array_29_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_6_clock),
    .reset(PE_Array_29_6_reset),
    .io_in_activate(PE_Array_29_6_io_in_activate),
    .io_in_weight(PE_Array_29_6_io_in_weight),
    .io_in_psum(PE_Array_29_6_io_in_psum),
    .io_in_flow(PE_Array_29_6_io_in_flow),
    .io_in_shift(PE_Array_29_6_io_in_shift),
    .io_out_activate(PE_Array_29_6_io_out_activate),
    .io_out_weight(PE_Array_29_6_io_out_weight),
    .io_out_psum(PE_Array_29_6_io_out_psum)
  );
  basic_PE PE_Array_29_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_7_clock),
    .reset(PE_Array_29_7_reset),
    .io_in_activate(PE_Array_29_7_io_in_activate),
    .io_in_weight(PE_Array_29_7_io_in_weight),
    .io_in_psum(PE_Array_29_7_io_in_psum),
    .io_in_flow(PE_Array_29_7_io_in_flow),
    .io_in_shift(PE_Array_29_7_io_in_shift),
    .io_out_activate(PE_Array_29_7_io_out_activate),
    .io_out_weight(PE_Array_29_7_io_out_weight),
    .io_out_psum(PE_Array_29_7_io_out_psum)
  );
  basic_PE PE_Array_29_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_8_clock),
    .reset(PE_Array_29_8_reset),
    .io_in_activate(PE_Array_29_8_io_in_activate),
    .io_in_weight(PE_Array_29_8_io_in_weight),
    .io_in_psum(PE_Array_29_8_io_in_psum),
    .io_in_flow(PE_Array_29_8_io_in_flow),
    .io_in_shift(PE_Array_29_8_io_in_shift),
    .io_out_activate(PE_Array_29_8_io_out_activate),
    .io_out_weight(PE_Array_29_8_io_out_weight),
    .io_out_psum(PE_Array_29_8_io_out_psum)
  );
  basic_PE PE_Array_29_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_9_clock),
    .reset(PE_Array_29_9_reset),
    .io_in_activate(PE_Array_29_9_io_in_activate),
    .io_in_weight(PE_Array_29_9_io_in_weight),
    .io_in_psum(PE_Array_29_9_io_in_psum),
    .io_in_flow(PE_Array_29_9_io_in_flow),
    .io_in_shift(PE_Array_29_9_io_in_shift),
    .io_out_activate(PE_Array_29_9_io_out_activate),
    .io_out_weight(PE_Array_29_9_io_out_weight),
    .io_out_psum(PE_Array_29_9_io_out_psum)
  );
  basic_PE PE_Array_29_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_10_clock),
    .reset(PE_Array_29_10_reset),
    .io_in_activate(PE_Array_29_10_io_in_activate),
    .io_in_weight(PE_Array_29_10_io_in_weight),
    .io_in_psum(PE_Array_29_10_io_in_psum),
    .io_in_flow(PE_Array_29_10_io_in_flow),
    .io_in_shift(PE_Array_29_10_io_in_shift),
    .io_out_activate(PE_Array_29_10_io_out_activate),
    .io_out_weight(PE_Array_29_10_io_out_weight),
    .io_out_psum(PE_Array_29_10_io_out_psum)
  );
  basic_PE PE_Array_29_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_11_clock),
    .reset(PE_Array_29_11_reset),
    .io_in_activate(PE_Array_29_11_io_in_activate),
    .io_in_weight(PE_Array_29_11_io_in_weight),
    .io_in_psum(PE_Array_29_11_io_in_psum),
    .io_in_flow(PE_Array_29_11_io_in_flow),
    .io_in_shift(PE_Array_29_11_io_in_shift),
    .io_out_activate(PE_Array_29_11_io_out_activate),
    .io_out_weight(PE_Array_29_11_io_out_weight),
    .io_out_psum(PE_Array_29_11_io_out_psum)
  );
  basic_PE PE_Array_29_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_12_clock),
    .reset(PE_Array_29_12_reset),
    .io_in_activate(PE_Array_29_12_io_in_activate),
    .io_in_weight(PE_Array_29_12_io_in_weight),
    .io_in_psum(PE_Array_29_12_io_in_psum),
    .io_in_flow(PE_Array_29_12_io_in_flow),
    .io_in_shift(PE_Array_29_12_io_in_shift),
    .io_out_activate(PE_Array_29_12_io_out_activate),
    .io_out_weight(PE_Array_29_12_io_out_weight),
    .io_out_psum(PE_Array_29_12_io_out_psum)
  );
  basic_PE PE_Array_29_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_13_clock),
    .reset(PE_Array_29_13_reset),
    .io_in_activate(PE_Array_29_13_io_in_activate),
    .io_in_weight(PE_Array_29_13_io_in_weight),
    .io_in_psum(PE_Array_29_13_io_in_psum),
    .io_in_flow(PE_Array_29_13_io_in_flow),
    .io_in_shift(PE_Array_29_13_io_in_shift),
    .io_out_activate(PE_Array_29_13_io_out_activate),
    .io_out_weight(PE_Array_29_13_io_out_weight),
    .io_out_psum(PE_Array_29_13_io_out_psum)
  );
  basic_PE PE_Array_29_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_14_clock),
    .reset(PE_Array_29_14_reset),
    .io_in_activate(PE_Array_29_14_io_in_activate),
    .io_in_weight(PE_Array_29_14_io_in_weight),
    .io_in_psum(PE_Array_29_14_io_in_psum),
    .io_in_flow(PE_Array_29_14_io_in_flow),
    .io_in_shift(PE_Array_29_14_io_in_shift),
    .io_out_activate(PE_Array_29_14_io_out_activate),
    .io_out_weight(PE_Array_29_14_io_out_weight),
    .io_out_psum(PE_Array_29_14_io_out_psum)
  );
  basic_PE PE_Array_29_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_15_clock),
    .reset(PE_Array_29_15_reset),
    .io_in_activate(PE_Array_29_15_io_in_activate),
    .io_in_weight(PE_Array_29_15_io_in_weight),
    .io_in_psum(PE_Array_29_15_io_in_psum),
    .io_in_flow(PE_Array_29_15_io_in_flow),
    .io_in_shift(PE_Array_29_15_io_in_shift),
    .io_out_activate(PE_Array_29_15_io_out_activate),
    .io_out_weight(PE_Array_29_15_io_out_weight),
    .io_out_psum(PE_Array_29_15_io_out_psum)
  );
  basic_PE PE_Array_29_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_16_clock),
    .reset(PE_Array_29_16_reset),
    .io_in_activate(PE_Array_29_16_io_in_activate),
    .io_in_weight(PE_Array_29_16_io_in_weight),
    .io_in_psum(PE_Array_29_16_io_in_psum),
    .io_in_flow(PE_Array_29_16_io_in_flow),
    .io_in_shift(PE_Array_29_16_io_in_shift),
    .io_out_activate(PE_Array_29_16_io_out_activate),
    .io_out_weight(PE_Array_29_16_io_out_weight),
    .io_out_psum(PE_Array_29_16_io_out_psum)
  );
  basic_PE PE_Array_29_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_17_clock),
    .reset(PE_Array_29_17_reset),
    .io_in_activate(PE_Array_29_17_io_in_activate),
    .io_in_weight(PE_Array_29_17_io_in_weight),
    .io_in_psum(PE_Array_29_17_io_in_psum),
    .io_in_flow(PE_Array_29_17_io_in_flow),
    .io_in_shift(PE_Array_29_17_io_in_shift),
    .io_out_activate(PE_Array_29_17_io_out_activate),
    .io_out_weight(PE_Array_29_17_io_out_weight),
    .io_out_psum(PE_Array_29_17_io_out_psum)
  );
  basic_PE PE_Array_29_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_18_clock),
    .reset(PE_Array_29_18_reset),
    .io_in_activate(PE_Array_29_18_io_in_activate),
    .io_in_weight(PE_Array_29_18_io_in_weight),
    .io_in_psum(PE_Array_29_18_io_in_psum),
    .io_in_flow(PE_Array_29_18_io_in_flow),
    .io_in_shift(PE_Array_29_18_io_in_shift),
    .io_out_activate(PE_Array_29_18_io_out_activate),
    .io_out_weight(PE_Array_29_18_io_out_weight),
    .io_out_psum(PE_Array_29_18_io_out_psum)
  );
  basic_PE PE_Array_29_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_19_clock),
    .reset(PE_Array_29_19_reset),
    .io_in_activate(PE_Array_29_19_io_in_activate),
    .io_in_weight(PE_Array_29_19_io_in_weight),
    .io_in_psum(PE_Array_29_19_io_in_psum),
    .io_in_flow(PE_Array_29_19_io_in_flow),
    .io_in_shift(PE_Array_29_19_io_in_shift),
    .io_out_activate(PE_Array_29_19_io_out_activate),
    .io_out_weight(PE_Array_29_19_io_out_weight),
    .io_out_psum(PE_Array_29_19_io_out_psum)
  );
  basic_PE PE_Array_29_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_20_clock),
    .reset(PE_Array_29_20_reset),
    .io_in_activate(PE_Array_29_20_io_in_activate),
    .io_in_weight(PE_Array_29_20_io_in_weight),
    .io_in_psum(PE_Array_29_20_io_in_psum),
    .io_in_flow(PE_Array_29_20_io_in_flow),
    .io_in_shift(PE_Array_29_20_io_in_shift),
    .io_out_activate(PE_Array_29_20_io_out_activate),
    .io_out_weight(PE_Array_29_20_io_out_weight),
    .io_out_psum(PE_Array_29_20_io_out_psum)
  );
  basic_PE PE_Array_29_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_21_clock),
    .reset(PE_Array_29_21_reset),
    .io_in_activate(PE_Array_29_21_io_in_activate),
    .io_in_weight(PE_Array_29_21_io_in_weight),
    .io_in_psum(PE_Array_29_21_io_in_psum),
    .io_in_flow(PE_Array_29_21_io_in_flow),
    .io_in_shift(PE_Array_29_21_io_in_shift),
    .io_out_activate(PE_Array_29_21_io_out_activate),
    .io_out_weight(PE_Array_29_21_io_out_weight),
    .io_out_psum(PE_Array_29_21_io_out_psum)
  );
  basic_PE PE_Array_29_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_22_clock),
    .reset(PE_Array_29_22_reset),
    .io_in_activate(PE_Array_29_22_io_in_activate),
    .io_in_weight(PE_Array_29_22_io_in_weight),
    .io_in_psum(PE_Array_29_22_io_in_psum),
    .io_in_flow(PE_Array_29_22_io_in_flow),
    .io_in_shift(PE_Array_29_22_io_in_shift),
    .io_out_activate(PE_Array_29_22_io_out_activate),
    .io_out_weight(PE_Array_29_22_io_out_weight),
    .io_out_psum(PE_Array_29_22_io_out_psum)
  );
  basic_PE PE_Array_29_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_23_clock),
    .reset(PE_Array_29_23_reset),
    .io_in_activate(PE_Array_29_23_io_in_activate),
    .io_in_weight(PE_Array_29_23_io_in_weight),
    .io_in_psum(PE_Array_29_23_io_in_psum),
    .io_in_flow(PE_Array_29_23_io_in_flow),
    .io_in_shift(PE_Array_29_23_io_in_shift),
    .io_out_activate(PE_Array_29_23_io_out_activate),
    .io_out_weight(PE_Array_29_23_io_out_weight),
    .io_out_psum(PE_Array_29_23_io_out_psum)
  );
  basic_PE PE_Array_29_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_24_clock),
    .reset(PE_Array_29_24_reset),
    .io_in_activate(PE_Array_29_24_io_in_activate),
    .io_in_weight(PE_Array_29_24_io_in_weight),
    .io_in_psum(PE_Array_29_24_io_in_psum),
    .io_in_flow(PE_Array_29_24_io_in_flow),
    .io_in_shift(PE_Array_29_24_io_in_shift),
    .io_out_activate(PE_Array_29_24_io_out_activate),
    .io_out_weight(PE_Array_29_24_io_out_weight),
    .io_out_psum(PE_Array_29_24_io_out_psum)
  );
  basic_PE PE_Array_29_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_25_clock),
    .reset(PE_Array_29_25_reset),
    .io_in_activate(PE_Array_29_25_io_in_activate),
    .io_in_weight(PE_Array_29_25_io_in_weight),
    .io_in_psum(PE_Array_29_25_io_in_psum),
    .io_in_flow(PE_Array_29_25_io_in_flow),
    .io_in_shift(PE_Array_29_25_io_in_shift),
    .io_out_activate(PE_Array_29_25_io_out_activate),
    .io_out_weight(PE_Array_29_25_io_out_weight),
    .io_out_psum(PE_Array_29_25_io_out_psum)
  );
  basic_PE PE_Array_29_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_26_clock),
    .reset(PE_Array_29_26_reset),
    .io_in_activate(PE_Array_29_26_io_in_activate),
    .io_in_weight(PE_Array_29_26_io_in_weight),
    .io_in_psum(PE_Array_29_26_io_in_psum),
    .io_in_flow(PE_Array_29_26_io_in_flow),
    .io_in_shift(PE_Array_29_26_io_in_shift),
    .io_out_activate(PE_Array_29_26_io_out_activate),
    .io_out_weight(PE_Array_29_26_io_out_weight),
    .io_out_psum(PE_Array_29_26_io_out_psum)
  );
  basic_PE PE_Array_29_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_27_clock),
    .reset(PE_Array_29_27_reset),
    .io_in_activate(PE_Array_29_27_io_in_activate),
    .io_in_weight(PE_Array_29_27_io_in_weight),
    .io_in_psum(PE_Array_29_27_io_in_psum),
    .io_in_flow(PE_Array_29_27_io_in_flow),
    .io_in_shift(PE_Array_29_27_io_in_shift),
    .io_out_activate(PE_Array_29_27_io_out_activate),
    .io_out_weight(PE_Array_29_27_io_out_weight),
    .io_out_psum(PE_Array_29_27_io_out_psum)
  );
  basic_PE PE_Array_29_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_28_clock),
    .reset(PE_Array_29_28_reset),
    .io_in_activate(PE_Array_29_28_io_in_activate),
    .io_in_weight(PE_Array_29_28_io_in_weight),
    .io_in_psum(PE_Array_29_28_io_in_psum),
    .io_in_flow(PE_Array_29_28_io_in_flow),
    .io_in_shift(PE_Array_29_28_io_in_shift),
    .io_out_activate(PE_Array_29_28_io_out_activate),
    .io_out_weight(PE_Array_29_28_io_out_weight),
    .io_out_psum(PE_Array_29_28_io_out_psum)
  );
  basic_PE PE_Array_29_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_29_clock),
    .reset(PE_Array_29_29_reset),
    .io_in_activate(PE_Array_29_29_io_in_activate),
    .io_in_weight(PE_Array_29_29_io_in_weight),
    .io_in_psum(PE_Array_29_29_io_in_psum),
    .io_in_flow(PE_Array_29_29_io_in_flow),
    .io_in_shift(PE_Array_29_29_io_in_shift),
    .io_out_activate(PE_Array_29_29_io_out_activate),
    .io_out_weight(PE_Array_29_29_io_out_weight),
    .io_out_psum(PE_Array_29_29_io_out_psum)
  );
  basic_PE PE_Array_29_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_30_clock),
    .reset(PE_Array_29_30_reset),
    .io_in_activate(PE_Array_29_30_io_in_activate),
    .io_in_weight(PE_Array_29_30_io_in_weight),
    .io_in_psum(PE_Array_29_30_io_in_psum),
    .io_in_flow(PE_Array_29_30_io_in_flow),
    .io_in_shift(PE_Array_29_30_io_in_shift),
    .io_out_activate(PE_Array_29_30_io_out_activate),
    .io_out_weight(PE_Array_29_30_io_out_weight),
    .io_out_psum(PE_Array_29_30_io_out_psum)
  );
  basic_PE PE_Array_29_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_29_31_clock),
    .reset(PE_Array_29_31_reset),
    .io_in_activate(PE_Array_29_31_io_in_activate),
    .io_in_weight(PE_Array_29_31_io_in_weight),
    .io_in_psum(PE_Array_29_31_io_in_psum),
    .io_in_flow(PE_Array_29_31_io_in_flow),
    .io_in_shift(PE_Array_29_31_io_in_shift),
    .io_out_activate(PE_Array_29_31_io_out_activate),
    .io_out_weight(PE_Array_29_31_io_out_weight),
    .io_out_psum(PE_Array_29_31_io_out_psum)
  );
  basic_PE PE_Array_30_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_0_clock),
    .reset(PE_Array_30_0_reset),
    .io_in_activate(PE_Array_30_0_io_in_activate),
    .io_in_weight(PE_Array_30_0_io_in_weight),
    .io_in_psum(PE_Array_30_0_io_in_psum),
    .io_in_flow(PE_Array_30_0_io_in_flow),
    .io_in_shift(PE_Array_30_0_io_in_shift),
    .io_out_activate(PE_Array_30_0_io_out_activate),
    .io_out_weight(PE_Array_30_0_io_out_weight),
    .io_out_psum(PE_Array_30_0_io_out_psum)
  );
  basic_PE PE_Array_30_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_1_clock),
    .reset(PE_Array_30_1_reset),
    .io_in_activate(PE_Array_30_1_io_in_activate),
    .io_in_weight(PE_Array_30_1_io_in_weight),
    .io_in_psum(PE_Array_30_1_io_in_psum),
    .io_in_flow(PE_Array_30_1_io_in_flow),
    .io_in_shift(PE_Array_30_1_io_in_shift),
    .io_out_activate(PE_Array_30_1_io_out_activate),
    .io_out_weight(PE_Array_30_1_io_out_weight),
    .io_out_psum(PE_Array_30_1_io_out_psum)
  );
  basic_PE PE_Array_30_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_2_clock),
    .reset(PE_Array_30_2_reset),
    .io_in_activate(PE_Array_30_2_io_in_activate),
    .io_in_weight(PE_Array_30_2_io_in_weight),
    .io_in_psum(PE_Array_30_2_io_in_psum),
    .io_in_flow(PE_Array_30_2_io_in_flow),
    .io_in_shift(PE_Array_30_2_io_in_shift),
    .io_out_activate(PE_Array_30_2_io_out_activate),
    .io_out_weight(PE_Array_30_2_io_out_weight),
    .io_out_psum(PE_Array_30_2_io_out_psum)
  );
  basic_PE PE_Array_30_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_3_clock),
    .reset(PE_Array_30_3_reset),
    .io_in_activate(PE_Array_30_3_io_in_activate),
    .io_in_weight(PE_Array_30_3_io_in_weight),
    .io_in_psum(PE_Array_30_3_io_in_psum),
    .io_in_flow(PE_Array_30_3_io_in_flow),
    .io_in_shift(PE_Array_30_3_io_in_shift),
    .io_out_activate(PE_Array_30_3_io_out_activate),
    .io_out_weight(PE_Array_30_3_io_out_weight),
    .io_out_psum(PE_Array_30_3_io_out_psum)
  );
  basic_PE PE_Array_30_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_4_clock),
    .reset(PE_Array_30_4_reset),
    .io_in_activate(PE_Array_30_4_io_in_activate),
    .io_in_weight(PE_Array_30_4_io_in_weight),
    .io_in_psum(PE_Array_30_4_io_in_psum),
    .io_in_flow(PE_Array_30_4_io_in_flow),
    .io_in_shift(PE_Array_30_4_io_in_shift),
    .io_out_activate(PE_Array_30_4_io_out_activate),
    .io_out_weight(PE_Array_30_4_io_out_weight),
    .io_out_psum(PE_Array_30_4_io_out_psum)
  );
  basic_PE PE_Array_30_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_5_clock),
    .reset(PE_Array_30_5_reset),
    .io_in_activate(PE_Array_30_5_io_in_activate),
    .io_in_weight(PE_Array_30_5_io_in_weight),
    .io_in_psum(PE_Array_30_5_io_in_psum),
    .io_in_flow(PE_Array_30_5_io_in_flow),
    .io_in_shift(PE_Array_30_5_io_in_shift),
    .io_out_activate(PE_Array_30_5_io_out_activate),
    .io_out_weight(PE_Array_30_5_io_out_weight),
    .io_out_psum(PE_Array_30_5_io_out_psum)
  );
  basic_PE PE_Array_30_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_6_clock),
    .reset(PE_Array_30_6_reset),
    .io_in_activate(PE_Array_30_6_io_in_activate),
    .io_in_weight(PE_Array_30_6_io_in_weight),
    .io_in_psum(PE_Array_30_6_io_in_psum),
    .io_in_flow(PE_Array_30_6_io_in_flow),
    .io_in_shift(PE_Array_30_6_io_in_shift),
    .io_out_activate(PE_Array_30_6_io_out_activate),
    .io_out_weight(PE_Array_30_6_io_out_weight),
    .io_out_psum(PE_Array_30_6_io_out_psum)
  );
  basic_PE PE_Array_30_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_7_clock),
    .reset(PE_Array_30_7_reset),
    .io_in_activate(PE_Array_30_7_io_in_activate),
    .io_in_weight(PE_Array_30_7_io_in_weight),
    .io_in_psum(PE_Array_30_7_io_in_psum),
    .io_in_flow(PE_Array_30_7_io_in_flow),
    .io_in_shift(PE_Array_30_7_io_in_shift),
    .io_out_activate(PE_Array_30_7_io_out_activate),
    .io_out_weight(PE_Array_30_7_io_out_weight),
    .io_out_psum(PE_Array_30_7_io_out_psum)
  );
  basic_PE PE_Array_30_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_8_clock),
    .reset(PE_Array_30_8_reset),
    .io_in_activate(PE_Array_30_8_io_in_activate),
    .io_in_weight(PE_Array_30_8_io_in_weight),
    .io_in_psum(PE_Array_30_8_io_in_psum),
    .io_in_flow(PE_Array_30_8_io_in_flow),
    .io_in_shift(PE_Array_30_8_io_in_shift),
    .io_out_activate(PE_Array_30_8_io_out_activate),
    .io_out_weight(PE_Array_30_8_io_out_weight),
    .io_out_psum(PE_Array_30_8_io_out_psum)
  );
  basic_PE PE_Array_30_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_9_clock),
    .reset(PE_Array_30_9_reset),
    .io_in_activate(PE_Array_30_9_io_in_activate),
    .io_in_weight(PE_Array_30_9_io_in_weight),
    .io_in_psum(PE_Array_30_9_io_in_psum),
    .io_in_flow(PE_Array_30_9_io_in_flow),
    .io_in_shift(PE_Array_30_9_io_in_shift),
    .io_out_activate(PE_Array_30_9_io_out_activate),
    .io_out_weight(PE_Array_30_9_io_out_weight),
    .io_out_psum(PE_Array_30_9_io_out_psum)
  );
  basic_PE PE_Array_30_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_10_clock),
    .reset(PE_Array_30_10_reset),
    .io_in_activate(PE_Array_30_10_io_in_activate),
    .io_in_weight(PE_Array_30_10_io_in_weight),
    .io_in_psum(PE_Array_30_10_io_in_psum),
    .io_in_flow(PE_Array_30_10_io_in_flow),
    .io_in_shift(PE_Array_30_10_io_in_shift),
    .io_out_activate(PE_Array_30_10_io_out_activate),
    .io_out_weight(PE_Array_30_10_io_out_weight),
    .io_out_psum(PE_Array_30_10_io_out_psum)
  );
  basic_PE PE_Array_30_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_11_clock),
    .reset(PE_Array_30_11_reset),
    .io_in_activate(PE_Array_30_11_io_in_activate),
    .io_in_weight(PE_Array_30_11_io_in_weight),
    .io_in_psum(PE_Array_30_11_io_in_psum),
    .io_in_flow(PE_Array_30_11_io_in_flow),
    .io_in_shift(PE_Array_30_11_io_in_shift),
    .io_out_activate(PE_Array_30_11_io_out_activate),
    .io_out_weight(PE_Array_30_11_io_out_weight),
    .io_out_psum(PE_Array_30_11_io_out_psum)
  );
  basic_PE PE_Array_30_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_12_clock),
    .reset(PE_Array_30_12_reset),
    .io_in_activate(PE_Array_30_12_io_in_activate),
    .io_in_weight(PE_Array_30_12_io_in_weight),
    .io_in_psum(PE_Array_30_12_io_in_psum),
    .io_in_flow(PE_Array_30_12_io_in_flow),
    .io_in_shift(PE_Array_30_12_io_in_shift),
    .io_out_activate(PE_Array_30_12_io_out_activate),
    .io_out_weight(PE_Array_30_12_io_out_weight),
    .io_out_psum(PE_Array_30_12_io_out_psum)
  );
  basic_PE PE_Array_30_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_13_clock),
    .reset(PE_Array_30_13_reset),
    .io_in_activate(PE_Array_30_13_io_in_activate),
    .io_in_weight(PE_Array_30_13_io_in_weight),
    .io_in_psum(PE_Array_30_13_io_in_psum),
    .io_in_flow(PE_Array_30_13_io_in_flow),
    .io_in_shift(PE_Array_30_13_io_in_shift),
    .io_out_activate(PE_Array_30_13_io_out_activate),
    .io_out_weight(PE_Array_30_13_io_out_weight),
    .io_out_psum(PE_Array_30_13_io_out_psum)
  );
  basic_PE PE_Array_30_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_14_clock),
    .reset(PE_Array_30_14_reset),
    .io_in_activate(PE_Array_30_14_io_in_activate),
    .io_in_weight(PE_Array_30_14_io_in_weight),
    .io_in_psum(PE_Array_30_14_io_in_psum),
    .io_in_flow(PE_Array_30_14_io_in_flow),
    .io_in_shift(PE_Array_30_14_io_in_shift),
    .io_out_activate(PE_Array_30_14_io_out_activate),
    .io_out_weight(PE_Array_30_14_io_out_weight),
    .io_out_psum(PE_Array_30_14_io_out_psum)
  );
  basic_PE PE_Array_30_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_15_clock),
    .reset(PE_Array_30_15_reset),
    .io_in_activate(PE_Array_30_15_io_in_activate),
    .io_in_weight(PE_Array_30_15_io_in_weight),
    .io_in_psum(PE_Array_30_15_io_in_psum),
    .io_in_flow(PE_Array_30_15_io_in_flow),
    .io_in_shift(PE_Array_30_15_io_in_shift),
    .io_out_activate(PE_Array_30_15_io_out_activate),
    .io_out_weight(PE_Array_30_15_io_out_weight),
    .io_out_psum(PE_Array_30_15_io_out_psum)
  );
  basic_PE PE_Array_30_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_16_clock),
    .reset(PE_Array_30_16_reset),
    .io_in_activate(PE_Array_30_16_io_in_activate),
    .io_in_weight(PE_Array_30_16_io_in_weight),
    .io_in_psum(PE_Array_30_16_io_in_psum),
    .io_in_flow(PE_Array_30_16_io_in_flow),
    .io_in_shift(PE_Array_30_16_io_in_shift),
    .io_out_activate(PE_Array_30_16_io_out_activate),
    .io_out_weight(PE_Array_30_16_io_out_weight),
    .io_out_psum(PE_Array_30_16_io_out_psum)
  );
  basic_PE PE_Array_30_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_17_clock),
    .reset(PE_Array_30_17_reset),
    .io_in_activate(PE_Array_30_17_io_in_activate),
    .io_in_weight(PE_Array_30_17_io_in_weight),
    .io_in_psum(PE_Array_30_17_io_in_psum),
    .io_in_flow(PE_Array_30_17_io_in_flow),
    .io_in_shift(PE_Array_30_17_io_in_shift),
    .io_out_activate(PE_Array_30_17_io_out_activate),
    .io_out_weight(PE_Array_30_17_io_out_weight),
    .io_out_psum(PE_Array_30_17_io_out_psum)
  );
  basic_PE PE_Array_30_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_18_clock),
    .reset(PE_Array_30_18_reset),
    .io_in_activate(PE_Array_30_18_io_in_activate),
    .io_in_weight(PE_Array_30_18_io_in_weight),
    .io_in_psum(PE_Array_30_18_io_in_psum),
    .io_in_flow(PE_Array_30_18_io_in_flow),
    .io_in_shift(PE_Array_30_18_io_in_shift),
    .io_out_activate(PE_Array_30_18_io_out_activate),
    .io_out_weight(PE_Array_30_18_io_out_weight),
    .io_out_psum(PE_Array_30_18_io_out_psum)
  );
  basic_PE PE_Array_30_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_19_clock),
    .reset(PE_Array_30_19_reset),
    .io_in_activate(PE_Array_30_19_io_in_activate),
    .io_in_weight(PE_Array_30_19_io_in_weight),
    .io_in_psum(PE_Array_30_19_io_in_psum),
    .io_in_flow(PE_Array_30_19_io_in_flow),
    .io_in_shift(PE_Array_30_19_io_in_shift),
    .io_out_activate(PE_Array_30_19_io_out_activate),
    .io_out_weight(PE_Array_30_19_io_out_weight),
    .io_out_psum(PE_Array_30_19_io_out_psum)
  );
  basic_PE PE_Array_30_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_20_clock),
    .reset(PE_Array_30_20_reset),
    .io_in_activate(PE_Array_30_20_io_in_activate),
    .io_in_weight(PE_Array_30_20_io_in_weight),
    .io_in_psum(PE_Array_30_20_io_in_psum),
    .io_in_flow(PE_Array_30_20_io_in_flow),
    .io_in_shift(PE_Array_30_20_io_in_shift),
    .io_out_activate(PE_Array_30_20_io_out_activate),
    .io_out_weight(PE_Array_30_20_io_out_weight),
    .io_out_psum(PE_Array_30_20_io_out_psum)
  );
  basic_PE PE_Array_30_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_21_clock),
    .reset(PE_Array_30_21_reset),
    .io_in_activate(PE_Array_30_21_io_in_activate),
    .io_in_weight(PE_Array_30_21_io_in_weight),
    .io_in_psum(PE_Array_30_21_io_in_psum),
    .io_in_flow(PE_Array_30_21_io_in_flow),
    .io_in_shift(PE_Array_30_21_io_in_shift),
    .io_out_activate(PE_Array_30_21_io_out_activate),
    .io_out_weight(PE_Array_30_21_io_out_weight),
    .io_out_psum(PE_Array_30_21_io_out_psum)
  );
  basic_PE PE_Array_30_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_22_clock),
    .reset(PE_Array_30_22_reset),
    .io_in_activate(PE_Array_30_22_io_in_activate),
    .io_in_weight(PE_Array_30_22_io_in_weight),
    .io_in_psum(PE_Array_30_22_io_in_psum),
    .io_in_flow(PE_Array_30_22_io_in_flow),
    .io_in_shift(PE_Array_30_22_io_in_shift),
    .io_out_activate(PE_Array_30_22_io_out_activate),
    .io_out_weight(PE_Array_30_22_io_out_weight),
    .io_out_psum(PE_Array_30_22_io_out_psum)
  );
  basic_PE PE_Array_30_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_23_clock),
    .reset(PE_Array_30_23_reset),
    .io_in_activate(PE_Array_30_23_io_in_activate),
    .io_in_weight(PE_Array_30_23_io_in_weight),
    .io_in_psum(PE_Array_30_23_io_in_psum),
    .io_in_flow(PE_Array_30_23_io_in_flow),
    .io_in_shift(PE_Array_30_23_io_in_shift),
    .io_out_activate(PE_Array_30_23_io_out_activate),
    .io_out_weight(PE_Array_30_23_io_out_weight),
    .io_out_psum(PE_Array_30_23_io_out_psum)
  );
  basic_PE PE_Array_30_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_24_clock),
    .reset(PE_Array_30_24_reset),
    .io_in_activate(PE_Array_30_24_io_in_activate),
    .io_in_weight(PE_Array_30_24_io_in_weight),
    .io_in_psum(PE_Array_30_24_io_in_psum),
    .io_in_flow(PE_Array_30_24_io_in_flow),
    .io_in_shift(PE_Array_30_24_io_in_shift),
    .io_out_activate(PE_Array_30_24_io_out_activate),
    .io_out_weight(PE_Array_30_24_io_out_weight),
    .io_out_psum(PE_Array_30_24_io_out_psum)
  );
  basic_PE PE_Array_30_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_25_clock),
    .reset(PE_Array_30_25_reset),
    .io_in_activate(PE_Array_30_25_io_in_activate),
    .io_in_weight(PE_Array_30_25_io_in_weight),
    .io_in_psum(PE_Array_30_25_io_in_psum),
    .io_in_flow(PE_Array_30_25_io_in_flow),
    .io_in_shift(PE_Array_30_25_io_in_shift),
    .io_out_activate(PE_Array_30_25_io_out_activate),
    .io_out_weight(PE_Array_30_25_io_out_weight),
    .io_out_psum(PE_Array_30_25_io_out_psum)
  );
  basic_PE PE_Array_30_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_26_clock),
    .reset(PE_Array_30_26_reset),
    .io_in_activate(PE_Array_30_26_io_in_activate),
    .io_in_weight(PE_Array_30_26_io_in_weight),
    .io_in_psum(PE_Array_30_26_io_in_psum),
    .io_in_flow(PE_Array_30_26_io_in_flow),
    .io_in_shift(PE_Array_30_26_io_in_shift),
    .io_out_activate(PE_Array_30_26_io_out_activate),
    .io_out_weight(PE_Array_30_26_io_out_weight),
    .io_out_psum(PE_Array_30_26_io_out_psum)
  );
  basic_PE PE_Array_30_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_27_clock),
    .reset(PE_Array_30_27_reset),
    .io_in_activate(PE_Array_30_27_io_in_activate),
    .io_in_weight(PE_Array_30_27_io_in_weight),
    .io_in_psum(PE_Array_30_27_io_in_psum),
    .io_in_flow(PE_Array_30_27_io_in_flow),
    .io_in_shift(PE_Array_30_27_io_in_shift),
    .io_out_activate(PE_Array_30_27_io_out_activate),
    .io_out_weight(PE_Array_30_27_io_out_weight),
    .io_out_psum(PE_Array_30_27_io_out_psum)
  );
  basic_PE PE_Array_30_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_28_clock),
    .reset(PE_Array_30_28_reset),
    .io_in_activate(PE_Array_30_28_io_in_activate),
    .io_in_weight(PE_Array_30_28_io_in_weight),
    .io_in_psum(PE_Array_30_28_io_in_psum),
    .io_in_flow(PE_Array_30_28_io_in_flow),
    .io_in_shift(PE_Array_30_28_io_in_shift),
    .io_out_activate(PE_Array_30_28_io_out_activate),
    .io_out_weight(PE_Array_30_28_io_out_weight),
    .io_out_psum(PE_Array_30_28_io_out_psum)
  );
  basic_PE PE_Array_30_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_29_clock),
    .reset(PE_Array_30_29_reset),
    .io_in_activate(PE_Array_30_29_io_in_activate),
    .io_in_weight(PE_Array_30_29_io_in_weight),
    .io_in_psum(PE_Array_30_29_io_in_psum),
    .io_in_flow(PE_Array_30_29_io_in_flow),
    .io_in_shift(PE_Array_30_29_io_in_shift),
    .io_out_activate(PE_Array_30_29_io_out_activate),
    .io_out_weight(PE_Array_30_29_io_out_weight),
    .io_out_psum(PE_Array_30_29_io_out_psum)
  );
  basic_PE PE_Array_30_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_30_clock),
    .reset(PE_Array_30_30_reset),
    .io_in_activate(PE_Array_30_30_io_in_activate),
    .io_in_weight(PE_Array_30_30_io_in_weight),
    .io_in_psum(PE_Array_30_30_io_in_psum),
    .io_in_flow(PE_Array_30_30_io_in_flow),
    .io_in_shift(PE_Array_30_30_io_in_shift),
    .io_out_activate(PE_Array_30_30_io_out_activate),
    .io_out_weight(PE_Array_30_30_io_out_weight),
    .io_out_psum(PE_Array_30_30_io_out_psum)
  );
  basic_PE PE_Array_30_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_30_31_clock),
    .reset(PE_Array_30_31_reset),
    .io_in_activate(PE_Array_30_31_io_in_activate),
    .io_in_weight(PE_Array_30_31_io_in_weight),
    .io_in_psum(PE_Array_30_31_io_in_psum),
    .io_in_flow(PE_Array_30_31_io_in_flow),
    .io_in_shift(PE_Array_30_31_io_in_shift),
    .io_out_activate(PE_Array_30_31_io_out_activate),
    .io_out_weight(PE_Array_30_31_io_out_weight),
    .io_out_psum(PE_Array_30_31_io_out_psum)
  );
  basic_PE PE_Array_31_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_0_clock),
    .reset(PE_Array_31_0_reset),
    .io_in_activate(PE_Array_31_0_io_in_activate),
    .io_in_weight(PE_Array_31_0_io_in_weight),
    .io_in_psum(PE_Array_31_0_io_in_psum),
    .io_in_flow(PE_Array_31_0_io_in_flow),
    .io_in_shift(PE_Array_31_0_io_in_shift),
    .io_out_activate(PE_Array_31_0_io_out_activate),
    .io_out_weight(PE_Array_31_0_io_out_weight),
    .io_out_psum(PE_Array_31_0_io_out_psum)
  );
  basic_PE PE_Array_31_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_1_clock),
    .reset(PE_Array_31_1_reset),
    .io_in_activate(PE_Array_31_1_io_in_activate),
    .io_in_weight(PE_Array_31_1_io_in_weight),
    .io_in_psum(PE_Array_31_1_io_in_psum),
    .io_in_flow(PE_Array_31_1_io_in_flow),
    .io_in_shift(PE_Array_31_1_io_in_shift),
    .io_out_activate(PE_Array_31_1_io_out_activate),
    .io_out_weight(PE_Array_31_1_io_out_weight),
    .io_out_psum(PE_Array_31_1_io_out_psum)
  );
  basic_PE PE_Array_31_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_2_clock),
    .reset(PE_Array_31_2_reset),
    .io_in_activate(PE_Array_31_2_io_in_activate),
    .io_in_weight(PE_Array_31_2_io_in_weight),
    .io_in_psum(PE_Array_31_2_io_in_psum),
    .io_in_flow(PE_Array_31_2_io_in_flow),
    .io_in_shift(PE_Array_31_2_io_in_shift),
    .io_out_activate(PE_Array_31_2_io_out_activate),
    .io_out_weight(PE_Array_31_2_io_out_weight),
    .io_out_psum(PE_Array_31_2_io_out_psum)
  );
  basic_PE PE_Array_31_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_3_clock),
    .reset(PE_Array_31_3_reset),
    .io_in_activate(PE_Array_31_3_io_in_activate),
    .io_in_weight(PE_Array_31_3_io_in_weight),
    .io_in_psum(PE_Array_31_3_io_in_psum),
    .io_in_flow(PE_Array_31_3_io_in_flow),
    .io_in_shift(PE_Array_31_3_io_in_shift),
    .io_out_activate(PE_Array_31_3_io_out_activate),
    .io_out_weight(PE_Array_31_3_io_out_weight),
    .io_out_psum(PE_Array_31_3_io_out_psum)
  );
  basic_PE PE_Array_31_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_4_clock),
    .reset(PE_Array_31_4_reset),
    .io_in_activate(PE_Array_31_4_io_in_activate),
    .io_in_weight(PE_Array_31_4_io_in_weight),
    .io_in_psum(PE_Array_31_4_io_in_psum),
    .io_in_flow(PE_Array_31_4_io_in_flow),
    .io_in_shift(PE_Array_31_4_io_in_shift),
    .io_out_activate(PE_Array_31_4_io_out_activate),
    .io_out_weight(PE_Array_31_4_io_out_weight),
    .io_out_psum(PE_Array_31_4_io_out_psum)
  );
  basic_PE PE_Array_31_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_5_clock),
    .reset(PE_Array_31_5_reset),
    .io_in_activate(PE_Array_31_5_io_in_activate),
    .io_in_weight(PE_Array_31_5_io_in_weight),
    .io_in_psum(PE_Array_31_5_io_in_psum),
    .io_in_flow(PE_Array_31_5_io_in_flow),
    .io_in_shift(PE_Array_31_5_io_in_shift),
    .io_out_activate(PE_Array_31_5_io_out_activate),
    .io_out_weight(PE_Array_31_5_io_out_weight),
    .io_out_psum(PE_Array_31_5_io_out_psum)
  );
  basic_PE PE_Array_31_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_6_clock),
    .reset(PE_Array_31_6_reset),
    .io_in_activate(PE_Array_31_6_io_in_activate),
    .io_in_weight(PE_Array_31_6_io_in_weight),
    .io_in_psum(PE_Array_31_6_io_in_psum),
    .io_in_flow(PE_Array_31_6_io_in_flow),
    .io_in_shift(PE_Array_31_6_io_in_shift),
    .io_out_activate(PE_Array_31_6_io_out_activate),
    .io_out_weight(PE_Array_31_6_io_out_weight),
    .io_out_psum(PE_Array_31_6_io_out_psum)
  );
  basic_PE PE_Array_31_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_7_clock),
    .reset(PE_Array_31_7_reset),
    .io_in_activate(PE_Array_31_7_io_in_activate),
    .io_in_weight(PE_Array_31_7_io_in_weight),
    .io_in_psum(PE_Array_31_7_io_in_psum),
    .io_in_flow(PE_Array_31_7_io_in_flow),
    .io_in_shift(PE_Array_31_7_io_in_shift),
    .io_out_activate(PE_Array_31_7_io_out_activate),
    .io_out_weight(PE_Array_31_7_io_out_weight),
    .io_out_psum(PE_Array_31_7_io_out_psum)
  );
  basic_PE PE_Array_31_8 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_8_clock),
    .reset(PE_Array_31_8_reset),
    .io_in_activate(PE_Array_31_8_io_in_activate),
    .io_in_weight(PE_Array_31_8_io_in_weight),
    .io_in_psum(PE_Array_31_8_io_in_psum),
    .io_in_flow(PE_Array_31_8_io_in_flow),
    .io_in_shift(PE_Array_31_8_io_in_shift),
    .io_out_activate(PE_Array_31_8_io_out_activate),
    .io_out_weight(PE_Array_31_8_io_out_weight),
    .io_out_psum(PE_Array_31_8_io_out_psum)
  );
  basic_PE PE_Array_31_9 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_9_clock),
    .reset(PE_Array_31_9_reset),
    .io_in_activate(PE_Array_31_9_io_in_activate),
    .io_in_weight(PE_Array_31_9_io_in_weight),
    .io_in_psum(PE_Array_31_9_io_in_psum),
    .io_in_flow(PE_Array_31_9_io_in_flow),
    .io_in_shift(PE_Array_31_9_io_in_shift),
    .io_out_activate(PE_Array_31_9_io_out_activate),
    .io_out_weight(PE_Array_31_9_io_out_weight),
    .io_out_psum(PE_Array_31_9_io_out_psum)
  );
  basic_PE PE_Array_31_10 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_10_clock),
    .reset(PE_Array_31_10_reset),
    .io_in_activate(PE_Array_31_10_io_in_activate),
    .io_in_weight(PE_Array_31_10_io_in_weight),
    .io_in_psum(PE_Array_31_10_io_in_psum),
    .io_in_flow(PE_Array_31_10_io_in_flow),
    .io_in_shift(PE_Array_31_10_io_in_shift),
    .io_out_activate(PE_Array_31_10_io_out_activate),
    .io_out_weight(PE_Array_31_10_io_out_weight),
    .io_out_psum(PE_Array_31_10_io_out_psum)
  );
  basic_PE PE_Array_31_11 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_11_clock),
    .reset(PE_Array_31_11_reset),
    .io_in_activate(PE_Array_31_11_io_in_activate),
    .io_in_weight(PE_Array_31_11_io_in_weight),
    .io_in_psum(PE_Array_31_11_io_in_psum),
    .io_in_flow(PE_Array_31_11_io_in_flow),
    .io_in_shift(PE_Array_31_11_io_in_shift),
    .io_out_activate(PE_Array_31_11_io_out_activate),
    .io_out_weight(PE_Array_31_11_io_out_weight),
    .io_out_psum(PE_Array_31_11_io_out_psum)
  );
  basic_PE PE_Array_31_12 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_12_clock),
    .reset(PE_Array_31_12_reset),
    .io_in_activate(PE_Array_31_12_io_in_activate),
    .io_in_weight(PE_Array_31_12_io_in_weight),
    .io_in_psum(PE_Array_31_12_io_in_psum),
    .io_in_flow(PE_Array_31_12_io_in_flow),
    .io_in_shift(PE_Array_31_12_io_in_shift),
    .io_out_activate(PE_Array_31_12_io_out_activate),
    .io_out_weight(PE_Array_31_12_io_out_weight),
    .io_out_psum(PE_Array_31_12_io_out_psum)
  );
  basic_PE PE_Array_31_13 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_13_clock),
    .reset(PE_Array_31_13_reset),
    .io_in_activate(PE_Array_31_13_io_in_activate),
    .io_in_weight(PE_Array_31_13_io_in_weight),
    .io_in_psum(PE_Array_31_13_io_in_psum),
    .io_in_flow(PE_Array_31_13_io_in_flow),
    .io_in_shift(PE_Array_31_13_io_in_shift),
    .io_out_activate(PE_Array_31_13_io_out_activate),
    .io_out_weight(PE_Array_31_13_io_out_weight),
    .io_out_psum(PE_Array_31_13_io_out_psum)
  );
  basic_PE PE_Array_31_14 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_14_clock),
    .reset(PE_Array_31_14_reset),
    .io_in_activate(PE_Array_31_14_io_in_activate),
    .io_in_weight(PE_Array_31_14_io_in_weight),
    .io_in_psum(PE_Array_31_14_io_in_psum),
    .io_in_flow(PE_Array_31_14_io_in_flow),
    .io_in_shift(PE_Array_31_14_io_in_shift),
    .io_out_activate(PE_Array_31_14_io_out_activate),
    .io_out_weight(PE_Array_31_14_io_out_weight),
    .io_out_psum(PE_Array_31_14_io_out_psum)
  );
  basic_PE PE_Array_31_15 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_15_clock),
    .reset(PE_Array_31_15_reset),
    .io_in_activate(PE_Array_31_15_io_in_activate),
    .io_in_weight(PE_Array_31_15_io_in_weight),
    .io_in_psum(PE_Array_31_15_io_in_psum),
    .io_in_flow(PE_Array_31_15_io_in_flow),
    .io_in_shift(PE_Array_31_15_io_in_shift),
    .io_out_activate(PE_Array_31_15_io_out_activate),
    .io_out_weight(PE_Array_31_15_io_out_weight),
    .io_out_psum(PE_Array_31_15_io_out_psum)
  );
  basic_PE PE_Array_31_16 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_16_clock),
    .reset(PE_Array_31_16_reset),
    .io_in_activate(PE_Array_31_16_io_in_activate),
    .io_in_weight(PE_Array_31_16_io_in_weight),
    .io_in_psum(PE_Array_31_16_io_in_psum),
    .io_in_flow(PE_Array_31_16_io_in_flow),
    .io_in_shift(PE_Array_31_16_io_in_shift),
    .io_out_activate(PE_Array_31_16_io_out_activate),
    .io_out_weight(PE_Array_31_16_io_out_weight),
    .io_out_psum(PE_Array_31_16_io_out_psum)
  );
  basic_PE PE_Array_31_17 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_17_clock),
    .reset(PE_Array_31_17_reset),
    .io_in_activate(PE_Array_31_17_io_in_activate),
    .io_in_weight(PE_Array_31_17_io_in_weight),
    .io_in_psum(PE_Array_31_17_io_in_psum),
    .io_in_flow(PE_Array_31_17_io_in_flow),
    .io_in_shift(PE_Array_31_17_io_in_shift),
    .io_out_activate(PE_Array_31_17_io_out_activate),
    .io_out_weight(PE_Array_31_17_io_out_weight),
    .io_out_psum(PE_Array_31_17_io_out_psum)
  );
  basic_PE PE_Array_31_18 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_18_clock),
    .reset(PE_Array_31_18_reset),
    .io_in_activate(PE_Array_31_18_io_in_activate),
    .io_in_weight(PE_Array_31_18_io_in_weight),
    .io_in_psum(PE_Array_31_18_io_in_psum),
    .io_in_flow(PE_Array_31_18_io_in_flow),
    .io_in_shift(PE_Array_31_18_io_in_shift),
    .io_out_activate(PE_Array_31_18_io_out_activate),
    .io_out_weight(PE_Array_31_18_io_out_weight),
    .io_out_psum(PE_Array_31_18_io_out_psum)
  );
  basic_PE PE_Array_31_19 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_19_clock),
    .reset(PE_Array_31_19_reset),
    .io_in_activate(PE_Array_31_19_io_in_activate),
    .io_in_weight(PE_Array_31_19_io_in_weight),
    .io_in_psum(PE_Array_31_19_io_in_psum),
    .io_in_flow(PE_Array_31_19_io_in_flow),
    .io_in_shift(PE_Array_31_19_io_in_shift),
    .io_out_activate(PE_Array_31_19_io_out_activate),
    .io_out_weight(PE_Array_31_19_io_out_weight),
    .io_out_psum(PE_Array_31_19_io_out_psum)
  );
  basic_PE PE_Array_31_20 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_20_clock),
    .reset(PE_Array_31_20_reset),
    .io_in_activate(PE_Array_31_20_io_in_activate),
    .io_in_weight(PE_Array_31_20_io_in_weight),
    .io_in_psum(PE_Array_31_20_io_in_psum),
    .io_in_flow(PE_Array_31_20_io_in_flow),
    .io_in_shift(PE_Array_31_20_io_in_shift),
    .io_out_activate(PE_Array_31_20_io_out_activate),
    .io_out_weight(PE_Array_31_20_io_out_weight),
    .io_out_psum(PE_Array_31_20_io_out_psum)
  );
  basic_PE PE_Array_31_21 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_21_clock),
    .reset(PE_Array_31_21_reset),
    .io_in_activate(PE_Array_31_21_io_in_activate),
    .io_in_weight(PE_Array_31_21_io_in_weight),
    .io_in_psum(PE_Array_31_21_io_in_psum),
    .io_in_flow(PE_Array_31_21_io_in_flow),
    .io_in_shift(PE_Array_31_21_io_in_shift),
    .io_out_activate(PE_Array_31_21_io_out_activate),
    .io_out_weight(PE_Array_31_21_io_out_weight),
    .io_out_psum(PE_Array_31_21_io_out_psum)
  );
  basic_PE PE_Array_31_22 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_22_clock),
    .reset(PE_Array_31_22_reset),
    .io_in_activate(PE_Array_31_22_io_in_activate),
    .io_in_weight(PE_Array_31_22_io_in_weight),
    .io_in_psum(PE_Array_31_22_io_in_psum),
    .io_in_flow(PE_Array_31_22_io_in_flow),
    .io_in_shift(PE_Array_31_22_io_in_shift),
    .io_out_activate(PE_Array_31_22_io_out_activate),
    .io_out_weight(PE_Array_31_22_io_out_weight),
    .io_out_psum(PE_Array_31_22_io_out_psum)
  );
  basic_PE PE_Array_31_23 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_23_clock),
    .reset(PE_Array_31_23_reset),
    .io_in_activate(PE_Array_31_23_io_in_activate),
    .io_in_weight(PE_Array_31_23_io_in_weight),
    .io_in_psum(PE_Array_31_23_io_in_psum),
    .io_in_flow(PE_Array_31_23_io_in_flow),
    .io_in_shift(PE_Array_31_23_io_in_shift),
    .io_out_activate(PE_Array_31_23_io_out_activate),
    .io_out_weight(PE_Array_31_23_io_out_weight),
    .io_out_psum(PE_Array_31_23_io_out_psum)
  );
  basic_PE PE_Array_31_24 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_24_clock),
    .reset(PE_Array_31_24_reset),
    .io_in_activate(PE_Array_31_24_io_in_activate),
    .io_in_weight(PE_Array_31_24_io_in_weight),
    .io_in_psum(PE_Array_31_24_io_in_psum),
    .io_in_flow(PE_Array_31_24_io_in_flow),
    .io_in_shift(PE_Array_31_24_io_in_shift),
    .io_out_activate(PE_Array_31_24_io_out_activate),
    .io_out_weight(PE_Array_31_24_io_out_weight),
    .io_out_psum(PE_Array_31_24_io_out_psum)
  );
  basic_PE PE_Array_31_25 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_25_clock),
    .reset(PE_Array_31_25_reset),
    .io_in_activate(PE_Array_31_25_io_in_activate),
    .io_in_weight(PE_Array_31_25_io_in_weight),
    .io_in_psum(PE_Array_31_25_io_in_psum),
    .io_in_flow(PE_Array_31_25_io_in_flow),
    .io_in_shift(PE_Array_31_25_io_in_shift),
    .io_out_activate(PE_Array_31_25_io_out_activate),
    .io_out_weight(PE_Array_31_25_io_out_weight),
    .io_out_psum(PE_Array_31_25_io_out_psum)
  );
  basic_PE PE_Array_31_26 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_26_clock),
    .reset(PE_Array_31_26_reset),
    .io_in_activate(PE_Array_31_26_io_in_activate),
    .io_in_weight(PE_Array_31_26_io_in_weight),
    .io_in_psum(PE_Array_31_26_io_in_psum),
    .io_in_flow(PE_Array_31_26_io_in_flow),
    .io_in_shift(PE_Array_31_26_io_in_shift),
    .io_out_activate(PE_Array_31_26_io_out_activate),
    .io_out_weight(PE_Array_31_26_io_out_weight),
    .io_out_psum(PE_Array_31_26_io_out_psum)
  );
  basic_PE PE_Array_31_27 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_27_clock),
    .reset(PE_Array_31_27_reset),
    .io_in_activate(PE_Array_31_27_io_in_activate),
    .io_in_weight(PE_Array_31_27_io_in_weight),
    .io_in_psum(PE_Array_31_27_io_in_psum),
    .io_in_flow(PE_Array_31_27_io_in_flow),
    .io_in_shift(PE_Array_31_27_io_in_shift),
    .io_out_activate(PE_Array_31_27_io_out_activate),
    .io_out_weight(PE_Array_31_27_io_out_weight),
    .io_out_psum(PE_Array_31_27_io_out_psum)
  );
  basic_PE PE_Array_31_28 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_28_clock),
    .reset(PE_Array_31_28_reset),
    .io_in_activate(PE_Array_31_28_io_in_activate),
    .io_in_weight(PE_Array_31_28_io_in_weight),
    .io_in_psum(PE_Array_31_28_io_in_psum),
    .io_in_flow(PE_Array_31_28_io_in_flow),
    .io_in_shift(PE_Array_31_28_io_in_shift),
    .io_out_activate(PE_Array_31_28_io_out_activate),
    .io_out_weight(PE_Array_31_28_io_out_weight),
    .io_out_psum(PE_Array_31_28_io_out_psum)
  );
  basic_PE PE_Array_31_29 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_29_clock),
    .reset(PE_Array_31_29_reset),
    .io_in_activate(PE_Array_31_29_io_in_activate),
    .io_in_weight(PE_Array_31_29_io_in_weight),
    .io_in_psum(PE_Array_31_29_io_in_psum),
    .io_in_flow(PE_Array_31_29_io_in_flow),
    .io_in_shift(PE_Array_31_29_io_in_shift),
    .io_out_activate(PE_Array_31_29_io_out_activate),
    .io_out_weight(PE_Array_31_29_io_out_weight),
    .io_out_psum(PE_Array_31_29_io_out_psum)
  );
  basic_PE PE_Array_31_30 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_30_clock),
    .reset(PE_Array_31_30_reset),
    .io_in_activate(PE_Array_31_30_io_in_activate),
    .io_in_weight(PE_Array_31_30_io_in_weight),
    .io_in_psum(PE_Array_31_30_io_in_psum),
    .io_in_flow(PE_Array_31_30_io_in_flow),
    .io_in_shift(PE_Array_31_30_io_in_shift),
    .io_out_activate(PE_Array_31_30_io_out_activate),
    .io_out_weight(PE_Array_31_30_io_out_weight),
    .io_out_psum(PE_Array_31_30_io_out_psum)
  );
  basic_PE PE_Array_31_31 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_31_31_clock),
    .reset(PE_Array_31_31_reset),
    .io_in_activate(PE_Array_31_31_io_in_activate),
    .io_in_weight(PE_Array_31_31_io_in_weight),
    .io_in_psum(PE_Array_31_31_io_in_psum),
    .io_in_flow(PE_Array_31_31_io_in_flow),
    .io_in_shift(PE_Array_31_31_io_in_shift),
    .io_out_activate(PE_Array_31_31_io_out_activate),
    .io_out_weight(PE_Array_31_31_io_out_weight),
    .io_out_psum(PE_Array_31_31_io_out_psum)
  );
  assign io_psum_0 = PE_Array_31_0_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_1 = PE_Array_31_1_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_2 = PE_Array_31_2_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_3 = PE_Array_31_3_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_4 = PE_Array_31_4_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_5 = PE_Array_31_5_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_6 = PE_Array_31_6_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_7 = PE_Array_31_7_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_8 = PE_Array_31_8_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_9 = PE_Array_31_9_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_10 = PE_Array_31_10_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_11 = PE_Array_31_11_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_12 = PE_Array_31_12_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_13 = PE_Array_31_13_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_14 = PE_Array_31_14_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_15 = PE_Array_31_15_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_16 = PE_Array_31_16_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_17 = PE_Array_31_17_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_18 = PE_Array_31_18_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_19 = PE_Array_31_19_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_20 = PE_Array_31_20_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_21 = PE_Array_31_21_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_22 = PE_Array_31_22_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_23 = PE_Array_31_23_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_24 = PE_Array_31_24_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_25 = PE_Array_31_25_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_26 = PE_Array_31_26_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_27 = PE_Array_31_27_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_28 = PE_Array_31_28_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_29 = PE_Array_31_29_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_30 = PE_Array_31_30_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_31 = PE_Array_31_31_io_out_psum; // @[DataPath.scala 24:10]
  assign io_valid_0 = valid_reg[0]; // @[Systolic_Array.scala 73:33]
  assign io_valid_1 = valid_reg[1]; // @[Systolic_Array.scala 73:33]
  assign io_valid_2 = valid_reg[2]; // @[Systolic_Array.scala 73:33]
  assign io_valid_3 = valid_reg[3]; // @[Systolic_Array.scala 73:33]
  assign io_valid_4 = valid_reg[4]; // @[Systolic_Array.scala 73:33]
  assign io_valid_5 = valid_reg[5]; // @[Systolic_Array.scala 73:33]
  assign io_valid_6 = valid_reg[6]; // @[Systolic_Array.scala 73:33]
  assign io_valid_7 = valid_reg[7]; // @[Systolic_Array.scala 73:33]
  assign io_valid_8 = valid_reg[8]; // @[Systolic_Array.scala 73:33]
  assign io_valid_9 = valid_reg[9]; // @[Systolic_Array.scala 73:33]
  assign io_valid_10 = valid_reg[10]; // @[Systolic_Array.scala 73:33]
  assign io_valid_11 = valid_reg[11]; // @[Systolic_Array.scala 73:33]
  assign io_valid_12 = valid_reg[12]; // @[Systolic_Array.scala 73:33]
  assign io_valid_13 = valid_reg[13]; // @[Systolic_Array.scala 73:33]
  assign io_valid_14 = valid_reg[14]; // @[Systolic_Array.scala 73:33]
  assign io_valid_15 = valid_reg[15]; // @[Systolic_Array.scala 73:33]
  assign io_valid_16 = valid_reg[16]; // @[Systolic_Array.scala 73:33]
  assign io_valid_17 = valid_reg[17]; // @[Systolic_Array.scala 73:33]
  assign io_valid_18 = valid_reg[18]; // @[Systolic_Array.scala 73:33]
  assign io_valid_19 = valid_reg[19]; // @[Systolic_Array.scala 73:33]
  assign io_valid_20 = valid_reg[20]; // @[Systolic_Array.scala 73:33]
  assign io_valid_21 = valid_reg[21]; // @[Systolic_Array.scala 73:33]
  assign io_valid_22 = valid_reg[22]; // @[Systolic_Array.scala 73:33]
  assign io_valid_23 = valid_reg[23]; // @[Systolic_Array.scala 73:33]
  assign io_valid_24 = valid_reg[24]; // @[Systolic_Array.scala 73:33]
  assign io_valid_25 = valid_reg[25]; // @[Systolic_Array.scala 73:33]
  assign io_valid_26 = valid_reg[26]; // @[Systolic_Array.scala 73:33]
  assign io_valid_27 = valid_reg[27]; // @[Systolic_Array.scala 73:33]
  assign io_valid_28 = valid_reg[28]; // @[Systolic_Array.scala 73:33]
  assign io_valid_29 = valid_reg[29]; // @[Systolic_Array.scala 73:33]
  assign io_valid_30 = valid_reg[30]; // @[Systolic_Array.scala 73:33]
  assign io_valid_31 = valid_reg[31]; // @[Systolic_Array.scala 73:33]
  assign PE_Array_0_0_clock = clock;
  assign PE_Array_0_0_reset = reset;
  assign PE_Array_0_0_io_in_activate = io_activate_0; // @[DataPath.scala 11:26]
  assign PE_Array_0_0_io_in_weight = io_weight_0; // @[DataPath.scala 20:23]
  assign PE_Array_0_0_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_1_clock = clock;
  assign PE_Array_0_1_reset = reset;
  assign PE_Array_0_1_io_in_activate = PE_Array_0_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_1_io_in_weight = io_weight_1; // @[DataPath.scala 20:23]
  assign PE_Array_0_1_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_2_clock = clock;
  assign PE_Array_0_2_reset = reset;
  assign PE_Array_0_2_io_in_activate = PE_Array_0_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_2_io_in_weight = io_weight_2; // @[DataPath.scala 20:23]
  assign PE_Array_0_2_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_3_clock = clock;
  assign PE_Array_0_3_reset = reset;
  assign PE_Array_0_3_io_in_activate = PE_Array_0_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_3_io_in_weight = io_weight_3; // @[DataPath.scala 20:23]
  assign PE_Array_0_3_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_4_clock = clock;
  assign PE_Array_0_4_reset = reset;
  assign PE_Array_0_4_io_in_activate = PE_Array_0_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_4_io_in_weight = io_weight_4; // @[DataPath.scala 20:23]
  assign PE_Array_0_4_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_5_clock = clock;
  assign PE_Array_0_5_reset = reset;
  assign PE_Array_0_5_io_in_activate = PE_Array_0_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_5_io_in_weight = io_weight_5; // @[DataPath.scala 20:23]
  assign PE_Array_0_5_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_6_clock = clock;
  assign PE_Array_0_6_reset = reset;
  assign PE_Array_0_6_io_in_activate = PE_Array_0_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_6_io_in_weight = io_weight_6; // @[DataPath.scala 20:23]
  assign PE_Array_0_6_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_7_clock = clock;
  assign PE_Array_0_7_reset = reset;
  assign PE_Array_0_7_io_in_activate = PE_Array_0_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_7_io_in_weight = io_weight_7; // @[DataPath.scala 20:23]
  assign PE_Array_0_7_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_8_clock = clock;
  assign PE_Array_0_8_reset = reset;
  assign PE_Array_0_8_io_in_activate = PE_Array_0_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_8_io_in_weight = io_weight_8; // @[DataPath.scala 20:23]
  assign PE_Array_0_8_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_9_clock = clock;
  assign PE_Array_0_9_reset = reset;
  assign PE_Array_0_9_io_in_activate = PE_Array_0_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_9_io_in_weight = io_weight_9; // @[DataPath.scala 20:23]
  assign PE_Array_0_9_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_10_clock = clock;
  assign PE_Array_0_10_reset = reset;
  assign PE_Array_0_10_io_in_activate = PE_Array_0_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_10_io_in_weight = io_weight_10; // @[DataPath.scala 20:23]
  assign PE_Array_0_10_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_11_clock = clock;
  assign PE_Array_0_11_reset = reset;
  assign PE_Array_0_11_io_in_activate = PE_Array_0_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_11_io_in_weight = io_weight_11; // @[DataPath.scala 20:23]
  assign PE_Array_0_11_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_12_clock = clock;
  assign PE_Array_0_12_reset = reset;
  assign PE_Array_0_12_io_in_activate = PE_Array_0_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_12_io_in_weight = io_weight_12; // @[DataPath.scala 20:23]
  assign PE_Array_0_12_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_13_clock = clock;
  assign PE_Array_0_13_reset = reset;
  assign PE_Array_0_13_io_in_activate = PE_Array_0_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_13_io_in_weight = io_weight_13; // @[DataPath.scala 20:23]
  assign PE_Array_0_13_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_14_clock = clock;
  assign PE_Array_0_14_reset = reset;
  assign PE_Array_0_14_io_in_activate = PE_Array_0_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_14_io_in_weight = io_weight_14; // @[DataPath.scala 20:23]
  assign PE_Array_0_14_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_15_clock = clock;
  assign PE_Array_0_15_reset = reset;
  assign PE_Array_0_15_io_in_activate = PE_Array_0_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_15_io_in_weight = io_weight_15; // @[DataPath.scala 20:23]
  assign PE_Array_0_15_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_16_clock = clock;
  assign PE_Array_0_16_reset = reset;
  assign PE_Array_0_16_io_in_activate = PE_Array_0_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_16_io_in_weight = io_weight_16; // @[DataPath.scala 20:23]
  assign PE_Array_0_16_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_17_clock = clock;
  assign PE_Array_0_17_reset = reset;
  assign PE_Array_0_17_io_in_activate = PE_Array_0_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_17_io_in_weight = io_weight_17; // @[DataPath.scala 20:23]
  assign PE_Array_0_17_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_18_clock = clock;
  assign PE_Array_0_18_reset = reset;
  assign PE_Array_0_18_io_in_activate = PE_Array_0_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_18_io_in_weight = io_weight_18; // @[DataPath.scala 20:23]
  assign PE_Array_0_18_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_19_clock = clock;
  assign PE_Array_0_19_reset = reset;
  assign PE_Array_0_19_io_in_activate = PE_Array_0_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_19_io_in_weight = io_weight_19; // @[DataPath.scala 20:23]
  assign PE_Array_0_19_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_20_clock = clock;
  assign PE_Array_0_20_reset = reset;
  assign PE_Array_0_20_io_in_activate = PE_Array_0_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_20_io_in_weight = io_weight_20; // @[DataPath.scala 20:23]
  assign PE_Array_0_20_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_21_clock = clock;
  assign PE_Array_0_21_reset = reset;
  assign PE_Array_0_21_io_in_activate = PE_Array_0_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_21_io_in_weight = io_weight_21; // @[DataPath.scala 20:23]
  assign PE_Array_0_21_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_22_clock = clock;
  assign PE_Array_0_22_reset = reset;
  assign PE_Array_0_22_io_in_activate = PE_Array_0_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_22_io_in_weight = io_weight_22; // @[DataPath.scala 20:23]
  assign PE_Array_0_22_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_23_clock = clock;
  assign PE_Array_0_23_reset = reset;
  assign PE_Array_0_23_io_in_activate = PE_Array_0_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_23_io_in_weight = io_weight_23; // @[DataPath.scala 20:23]
  assign PE_Array_0_23_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_24_clock = clock;
  assign PE_Array_0_24_reset = reset;
  assign PE_Array_0_24_io_in_activate = PE_Array_0_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_24_io_in_weight = io_weight_24; // @[DataPath.scala 20:23]
  assign PE_Array_0_24_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_25_clock = clock;
  assign PE_Array_0_25_reset = reset;
  assign PE_Array_0_25_io_in_activate = PE_Array_0_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_25_io_in_weight = io_weight_25; // @[DataPath.scala 20:23]
  assign PE_Array_0_25_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_26_clock = clock;
  assign PE_Array_0_26_reset = reset;
  assign PE_Array_0_26_io_in_activate = PE_Array_0_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_26_io_in_weight = io_weight_26; // @[DataPath.scala 20:23]
  assign PE_Array_0_26_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_27_clock = clock;
  assign PE_Array_0_27_reset = reset;
  assign PE_Array_0_27_io_in_activate = PE_Array_0_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_27_io_in_weight = io_weight_27; // @[DataPath.scala 20:23]
  assign PE_Array_0_27_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_28_clock = clock;
  assign PE_Array_0_28_reset = reset;
  assign PE_Array_0_28_io_in_activate = PE_Array_0_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_28_io_in_weight = io_weight_28; // @[DataPath.scala 20:23]
  assign PE_Array_0_28_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_29_clock = clock;
  assign PE_Array_0_29_reset = reset;
  assign PE_Array_0_29_io_in_activate = PE_Array_0_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_29_io_in_weight = io_weight_29; // @[DataPath.scala 20:23]
  assign PE_Array_0_29_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_30_clock = clock;
  assign PE_Array_0_30_reset = reset;
  assign PE_Array_0_30_io_in_activate = PE_Array_0_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_30_io_in_weight = io_weight_30; // @[DataPath.scala 20:23]
  assign PE_Array_0_30_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_31_clock = clock;
  assign PE_Array_0_31_reset = reset;
  assign PE_Array_0_31_io_in_activate = PE_Array_0_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_31_io_in_weight = io_weight_31; // @[DataPath.scala 20:23]
  assign PE_Array_0_31_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_0_clock = clock;
  assign PE_Array_1_0_reset = reset;
  assign PE_Array_1_0_io_in_activate = io_activate_1; // @[DataPath.scala 11:26]
  assign PE_Array_1_0_io_in_weight = PE_Array_0_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_0_io_in_psum = PE_Array_0_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_1_clock = clock;
  assign PE_Array_1_1_reset = reset;
  assign PE_Array_1_1_io_in_activate = PE_Array_1_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_1_io_in_weight = PE_Array_0_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_1_io_in_psum = PE_Array_0_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_2_clock = clock;
  assign PE_Array_1_2_reset = reset;
  assign PE_Array_1_2_io_in_activate = PE_Array_1_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_2_io_in_weight = PE_Array_0_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_2_io_in_psum = PE_Array_0_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_3_clock = clock;
  assign PE_Array_1_3_reset = reset;
  assign PE_Array_1_3_io_in_activate = PE_Array_1_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_3_io_in_weight = PE_Array_0_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_3_io_in_psum = PE_Array_0_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_4_clock = clock;
  assign PE_Array_1_4_reset = reset;
  assign PE_Array_1_4_io_in_activate = PE_Array_1_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_4_io_in_weight = PE_Array_0_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_4_io_in_psum = PE_Array_0_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_5_clock = clock;
  assign PE_Array_1_5_reset = reset;
  assign PE_Array_1_5_io_in_activate = PE_Array_1_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_5_io_in_weight = PE_Array_0_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_5_io_in_psum = PE_Array_0_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_6_clock = clock;
  assign PE_Array_1_6_reset = reset;
  assign PE_Array_1_6_io_in_activate = PE_Array_1_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_6_io_in_weight = PE_Array_0_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_6_io_in_psum = PE_Array_0_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_7_clock = clock;
  assign PE_Array_1_7_reset = reset;
  assign PE_Array_1_7_io_in_activate = PE_Array_1_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_7_io_in_weight = PE_Array_0_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_7_io_in_psum = PE_Array_0_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_8_clock = clock;
  assign PE_Array_1_8_reset = reset;
  assign PE_Array_1_8_io_in_activate = PE_Array_1_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_8_io_in_weight = PE_Array_0_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_8_io_in_psum = PE_Array_0_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_9_clock = clock;
  assign PE_Array_1_9_reset = reset;
  assign PE_Array_1_9_io_in_activate = PE_Array_1_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_9_io_in_weight = PE_Array_0_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_9_io_in_psum = PE_Array_0_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_10_clock = clock;
  assign PE_Array_1_10_reset = reset;
  assign PE_Array_1_10_io_in_activate = PE_Array_1_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_10_io_in_weight = PE_Array_0_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_10_io_in_psum = PE_Array_0_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_11_clock = clock;
  assign PE_Array_1_11_reset = reset;
  assign PE_Array_1_11_io_in_activate = PE_Array_1_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_11_io_in_weight = PE_Array_0_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_11_io_in_psum = PE_Array_0_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_12_clock = clock;
  assign PE_Array_1_12_reset = reset;
  assign PE_Array_1_12_io_in_activate = PE_Array_1_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_12_io_in_weight = PE_Array_0_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_12_io_in_psum = PE_Array_0_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_13_clock = clock;
  assign PE_Array_1_13_reset = reset;
  assign PE_Array_1_13_io_in_activate = PE_Array_1_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_13_io_in_weight = PE_Array_0_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_13_io_in_psum = PE_Array_0_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_14_clock = clock;
  assign PE_Array_1_14_reset = reset;
  assign PE_Array_1_14_io_in_activate = PE_Array_1_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_14_io_in_weight = PE_Array_0_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_14_io_in_psum = PE_Array_0_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_15_clock = clock;
  assign PE_Array_1_15_reset = reset;
  assign PE_Array_1_15_io_in_activate = PE_Array_1_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_15_io_in_weight = PE_Array_0_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_15_io_in_psum = PE_Array_0_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_16_clock = clock;
  assign PE_Array_1_16_reset = reset;
  assign PE_Array_1_16_io_in_activate = PE_Array_1_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_16_io_in_weight = PE_Array_0_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_16_io_in_psum = PE_Array_0_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_17_clock = clock;
  assign PE_Array_1_17_reset = reset;
  assign PE_Array_1_17_io_in_activate = PE_Array_1_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_17_io_in_weight = PE_Array_0_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_17_io_in_psum = PE_Array_0_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_18_clock = clock;
  assign PE_Array_1_18_reset = reset;
  assign PE_Array_1_18_io_in_activate = PE_Array_1_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_18_io_in_weight = PE_Array_0_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_18_io_in_psum = PE_Array_0_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_19_clock = clock;
  assign PE_Array_1_19_reset = reset;
  assign PE_Array_1_19_io_in_activate = PE_Array_1_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_19_io_in_weight = PE_Array_0_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_19_io_in_psum = PE_Array_0_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_20_clock = clock;
  assign PE_Array_1_20_reset = reset;
  assign PE_Array_1_20_io_in_activate = PE_Array_1_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_20_io_in_weight = PE_Array_0_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_20_io_in_psum = PE_Array_0_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_21_clock = clock;
  assign PE_Array_1_21_reset = reset;
  assign PE_Array_1_21_io_in_activate = PE_Array_1_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_21_io_in_weight = PE_Array_0_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_21_io_in_psum = PE_Array_0_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_22_clock = clock;
  assign PE_Array_1_22_reset = reset;
  assign PE_Array_1_22_io_in_activate = PE_Array_1_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_22_io_in_weight = PE_Array_0_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_22_io_in_psum = PE_Array_0_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_23_clock = clock;
  assign PE_Array_1_23_reset = reset;
  assign PE_Array_1_23_io_in_activate = PE_Array_1_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_23_io_in_weight = PE_Array_0_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_23_io_in_psum = PE_Array_0_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_24_clock = clock;
  assign PE_Array_1_24_reset = reset;
  assign PE_Array_1_24_io_in_activate = PE_Array_1_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_24_io_in_weight = PE_Array_0_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_24_io_in_psum = PE_Array_0_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_25_clock = clock;
  assign PE_Array_1_25_reset = reset;
  assign PE_Array_1_25_io_in_activate = PE_Array_1_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_25_io_in_weight = PE_Array_0_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_25_io_in_psum = PE_Array_0_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_26_clock = clock;
  assign PE_Array_1_26_reset = reset;
  assign PE_Array_1_26_io_in_activate = PE_Array_1_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_26_io_in_weight = PE_Array_0_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_26_io_in_psum = PE_Array_0_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_27_clock = clock;
  assign PE_Array_1_27_reset = reset;
  assign PE_Array_1_27_io_in_activate = PE_Array_1_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_27_io_in_weight = PE_Array_0_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_27_io_in_psum = PE_Array_0_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_28_clock = clock;
  assign PE_Array_1_28_reset = reset;
  assign PE_Array_1_28_io_in_activate = PE_Array_1_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_28_io_in_weight = PE_Array_0_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_28_io_in_psum = PE_Array_0_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_29_clock = clock;
  assign PE_Array_1_29_reset = reset;
  assign PE_Array_1_29_io_in_activate = PE_Array_1_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_29_io_in_weight = PE_Array_0_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_29_io_in_psum = PE_Array_0_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_30_clock = clock;
  assign PE_Array_1_30_reset = reset;
  assign PE_Array_1_30_io_in_activate = PE_Array_1_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_30_io_in_weight = PE_Array_0_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_30_io_in_psum = PE_Array_0_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_31_clock = clock;
  assign PE_Array_1_31_reset = reset;
  assign PE_Array_1_31_io_in_activate = PE_Array_1_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_31_io_in_weight = PE_Array_0_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_31_io_in_psum = PE_Array_0_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_0_clock = clock;
  assign PE_Array_2_0_reset = reset;
  assign PE_Array_2_0_io_in_activate = io_activate_2; // @[DataPath.scala 11:26]
  assign PE_Array_2_0_io_in_weight = PE_Array_1_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_0_io_in_psum = PE_Array_1_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_1_clock = clock;
  assign PE_Array_2_1_reset = reset;
  assign PE_Array_2_1_io_in_activate = PE_Array_2_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_1_io_in_weight = PE_Array_1_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_1_io_in_psum = PE_Array_1_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_2_clock = clock;
  assign PE_Array_2_2_reset = reset;
  assign PE_Array_2_2_io_in_activate = PE_Array_2_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_2_io_in_weight = PE_Array_1_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_2_io_in_psum = PE_Array_1_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_3_clock = clock;
  assign PE_Array_2_3_reset = reset;
  assign PE_Array_2_3_io_in_activate = PE_Array_2_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_3_io_in_weight = PE_Array_1_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_3_io_in_psum = PE_Array_1_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_4_clock = clock;
  assign PE_Array_2_4_reset = reset;
  assign PE_Array_2_4_io_in_activate = PE_Array_2_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_4_io_in_weight = PE_Array_1_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_4_io_in_psum = PE_Array_1_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_5_clock = clock;
  assign PE_Array_2_5_reset = reset;
  assign PE_Array_2_5_io_in_activate = PE_Array_2_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_5_io_in_weight = PE_Array_1_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_5_io_in_psum = PE_Array_1_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_6_clock = clock;
  assign PE_Array_2_6_reset = reset;
  assign PE_Array_2_6_io_in_activate = PE_Array_2_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_6_io_in_weight = PE_Array_1_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_6_io_in_psum = PE_Array_1_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_7_clock = clock;
  assign PE_Array_2_7_reset = reset;
  assign PE_Array_2_7_io_in_activate = PE_Array_2_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_7_io_in_weight = PE_Array_1_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_7_io_in_psum = PE_Array_1_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_8_clock = clock;
  assign PE_Array_2_8_reset = reset;
  assign PE_Array_2_8_io_in_activate = PE_Array_2_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_8_io_in_weight = PE_Array_1_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_8_io_in_psum = PE_Array_1_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_9_clock = clock;
  assign PE_Array_2_9_reset = reset;
  assign PE_Array_2_9_io_in_activate = PE_Array_2_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_9_io_in_weight = PE_Array_1_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_9_io_in_psum = PE_Array_1_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_10_clock = clock;
  assign PE_Array_2_10_reset = reset;
  assign PE_Array_2_10_io_in_activate = PE_Array_2_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_10_io_in_weight = PE_Array_1_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_10_io_in_psum = PE_Array_1_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_11_clock = clock;
  assign PE_Array_2_11_reset = reset;
  assign PE_Array_2_11_io_in_activate = PE_Array_2_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_11_io_in_weight = PE_Array_1_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_11_io_in_psum = PE_Array_1_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_12_clock = clock;
  assign PE_Array_2_12_reset = reset;
  assign PE_Array_2_12_io_in_activate = PE_Array_2_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_12_io_in_weight = PE_Array_1_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_12_io_in_psum = PE_Array_1_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_13_clock = clock;
  assign PE_Array_2_13_reset = reset;
  assign PE_Array_2_13_io_in_activate = PE_Array_2_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_13_io_in_weight = PE_Array_1_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_13_io_in_psum = PE_Array_1_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_14_clock = clock;
  assign PE_Array_2_14_reset = reset;
  assign PE_Array_2_14_io_in_activate = PE_Array_2_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_14_io_in_weight = PE_Array_1_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_14_io_in_psum = PE_Array_1_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_15_clock = clock;
  assign PE_Array_2_15_reset = reset;
  assign PE_Array_2_15_io_in_activate = PE_Array_2_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_15_io_in_weight = PE_Array_1_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_15_io_in_psum = PE_Array_1_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_16_clock = clock;
  assign PE_Array_2_16_reset = reset;
  assign PE_Array_2_16_io_in_activate = PE_Array_2_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_16_io_in_weight = PE_Array_1_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_16_io_in_psum = PE_Array_1_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_17_clock = clock;
  assign PE_Array_2_17_reset = reset;
  assign PE_Array_2_17_io_in_activate = PE_Array_2_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_17_io_in_weight = PE_Array_1_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_17_io_in_psum = PE_Array_1_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_18_clock = clock;
  assign PE_Array_2_18_reset = reset;
  assign PE_Array_2_18_io_in_activate = PE_Array_2_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_18_io_in_weight = PE_Array_1_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_18_io_in_psum = PE_Array_1_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_19_clock = clock;
  assign PE_Array_2_19_reset = reset;
  assign PE_Array_2_19_io_in_activate = PE_Array_2_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_19_io_in_weight = PE_Array_1_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_19_io_in_psum = PE_Array_1_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_20_clock = clock;
  assign PE_Array_2_20_reset = reset;
  assign PE_Array_2_20_io_in_activate = PE_Array_2_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_20_io_in_weight = PE_Array_1_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_20_io_in_psum = PE_Array_1_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_21_clock = clock;
  assign PE_Array_2_21_reset = reset;
  assign PE_Array_2_21_io_in_activate = PE_Array_2_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_21_io_in_weight = PE_Array_1_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_21_io_in_psum = PE_Array_1_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_22_clock = clock;
  assign PE_Array_2_22_reset = reset;
  assign PE_Array_2_22_io_in_activate = PE_Array_2_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_22_io_in_weight = PE_Array_1_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_22_io_in_psum = PE_Array_1_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_23_clock = clock;
  assign PE_Array_2_23_reset = reset;
  assign PE_Array_2_23_io_in_activate = PE_Array_2_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_23_io_in_weight = PE_Array_1_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_23_io_in_psum = PE_Array_1_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_24_clock = clock;
  assign PE_Array_2_24_reset = reset;
  assign PE_Array_2_24_io_in_activate = PE_Array_2_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_24_io_in_weight = PE_Array_1_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_24_io_in_psum = PE_Array_1_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_25_clock = clock;
  assign PE_Array_2_25_reset = reset;
  assign PE_Array_2_25_io_in_activate = PE_Array_2_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_25_io_in_weight = PE_Array_1_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_25_io_in_psum = PE_Array_1_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_26_clock = clock;
  assign PE_Array_2_26_reset = reset;
  assign PE_Array_2_26_io_in_activate = PE_Array_2_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_26_io_in_weight = PE_Array_1_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_26_io_in_psum = PE_Array_1_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_27_clock = clock;
  assign PE_Array_2_27_reset = reset;
  assign PE_Array_2_27_io_in_activate = PE_Array_2_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_27_io_in_weight = PE_Array_1_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_27_io_in_psum = PE_Array_1_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_28_clock = clock;
  assign PE_Array_2_28_reset = reset;
  assign PE_Array_2_28_io_in_activate = PE_Array_2_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_28_io_in_weight = PE_Array_1_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_28_io_in_psum = PE_Array_1_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_29_clock = clock;
  assign PE_Array_2_29_reset = reset;
  assign PE_Array_2_29_io_in_activate = PE_Array_2_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_29_io_in_weight = PE_Array_1_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_29_io_in_psum = PE_Array_1_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_30_clock = clock;
  assign PE_Array_2_30_reset = reset;
  assign PE_Array_2_30_io_in_activate = PE_Array_2_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_30_io_in_weight = PE_Array_1_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_30_io_in_psum = PE_Array_1_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_31_clock = clock;
  assign PE_Array_2_31_reset = reset;
  assign PE_Array_2_31_io_in_activate = PE_Array_2_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_31_io_in_weight = PE_Array_1_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_31_io_in_psum = PE_Array_1_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_0_clock = clock;
  assign PE_Array_3_0_reset = reset;
  assign PE_Array_3_0_io_in_activate = io_activate_3; // @[DataPath.scala 11:26]
  assign PE_Array_3_0_io_in_weight = PE_Array_2_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_0_io_in_psum = PE_Array_2_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_1_clock = clock;
  assign PE_Array_3_1_reset = reset;
  assign PE_Array_3_1_io_in_activate = PE_Array_3_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_1_io_in_weight = PE_Array_2_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_1_io_in_psum = PE_Array_2_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_2_clock = clock;
  assign PE_Array_3_2_reset = reset;
  assign PE_Array_3_2_io_in_activate = PE_Array_3_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_2_io_in_weight = PE_Array_2_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_2_io_in_psum = PE_Array_2_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_3_clock = clock;
  assign PE_Array_3_3_reset = reset;
  assign PE_Array_3_3_io_in_activate = PE_Array_3_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_3_io_in_weight = PE_Array_2_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_3_io_in_psum = PE_Array_2_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_4_clock = clock;
  assign PE_Array_3_4_reset = reset;
  assign PE_Array_3_4_io_in_activate = PE_Array_3_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_4_io_in_weight = PE_Array_2_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_4_io_in_psum = PE_Array_2_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_5_clock = clock;
  assign PE_Array_3_5_reset = reset;
  assign PE_Array_3_5_io_in_activate = PE_Array_3_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_5_io_in_weight = PE_Array_2_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_5_io_in_psum = PE_Array_2_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_6_clock = clock;
  assign PE_Array_3_6_reset = reset;
  assign PE_Array_3_6_io_in_activate = PE_Array_3_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_6_io_in_weight = PE_Array_2_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_6_io_in_psum = PE_Array_2_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_7_clock = clock;
  assign PE_Array_3_7_reset = reset;
  assign PE_Array_3_7_io_in_activate = PE_Array_3_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_7_io_in_weight = PE_Array_2_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_7_io_in_psum = PE_Array_2_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_8_clock = clock;
  assign PE_Array_3_8_reset = reset;
  assign PE_Array_3_8_io_in_activate = PE_Array_3_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_8_io_in_weight = PE_Array_2_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_8_io_in_psum = PE_Array_2_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_9_clock = clock;
  assign PE_Array_3_9_reset = reset;
  assign PE_Array_3_9_io_in_activate = PE_Array_3_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_9_io_in_weight = PE_Array_2_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_9_io_in_psum = PE_Array_2_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_10_clock = clock;
  assign PE_Array_3_10_reset = reset;
  assign PE_Array_3_10_io_in_activate = PE_Array_3_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_10_io_in_weight = PE_Array_2_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_10_io_in_psum = PE_Array_2_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_11_clock = clock;
  assign PE_Array_3_11_reset = reset;
  assign PE_Array_3_11_io_in_activate = PE_Array_3_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_11_io_in_weight = PE_Array_2_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_11_io_in_psum = PE_Array_2_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_12_clock = clock;
  assign PE_Array_3_12_reset = reset;
  assign PE_Array_3_12_io_in_activate = PE_Array_3_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_12_io_in_weight = PE_Array_2_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_12_io_in_psum = PE_Array_2_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_13_clock = clock;
  assign PE_Array_3_13_reset = reset;
  assign PE_Array_3_13_io_in_activate = PE_Array_3_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_13_io_in_weight = PE_Array_2_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_13_io_in_psum = PE_Array_2_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_14_clock = clock;
  assign PE_Array_3_14_reset = reset;
  assign PE_Array_3_14_io_in_activate = PE_Array_3_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_14_io_in_weight = PE_Array_2_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_14_io_in_psum = PE_Array_2_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_15_clock = clock;
  assign PE_Array_3_15_reset = reset;
  assign PE_Array_3_15_io_in_activate = PE_Array_3_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_15_io_in_weight = PE_Array_2_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_15_io_in_psum = PE_Array_2_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_16_clock = clock;
  assign PE_Array_3_16_reset = reset;
  assign PE_Array_3_16_io_in_activate = PE_Array_3_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_16_io_in_weight = PE_Array_2_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_16_io_in_psum = PE_Array_2_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_17_clock = clock;
  assign PE_Array_3_17_reset = reset;
  assign PE_Array_3_17_io_in_activate = PE_Array_3_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_17_io_in_weight = PE_Array_2_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_17_io_in_psum = PE_Array_2_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_18_clock = clock;
  assign PE_Array_3_18_reset = reset;
  assign PE_Array_3_18_io_in_activate = PE_Array_3_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_18_io_in_weight = PE_Array_2_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_18_io_in_psum = PE_Array_2_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_19_clock = clock;
  assign PE_Array_3_19_reset = reset;
  assign PE_Array_3_19_io_in_activate = PE_Array_3_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_19_io_in_weight = PE_Array_2_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_19_io_in_psum = PE_Array_2_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_20_clock = clock;
  assign PE_Array_3_20_reset = reset;
  assign PE_Array_3_20_io_in_activate = PE_Array_3_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_20_io_in_weight = PE_Array_2_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_20_io_in_psum = PE_Array_2_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_21_clock = clock;
  assign PE_Array_3_21_reset = reset;
  assign PE_Array_3_21_io_in_activate = PE_Array_3_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_21_io_in_weight = PE_Array_2_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_21_io_in_psum = PE_Array_2_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_22_clock = clock;
  assign PE_Array_3_22_reset = reset;
  assign PE_Array_3_22_io_in_activate = PE_Array_3_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_22_io_in_weight = PE_Array_2_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_22_io_in_psum = PE_Array_2_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_23_clock = clock;
  assign PE_Array_3_23_reset = reset;
  assign PE_Array_3_23_io_in_activate = PE_Array_3_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_23_io_in_weight = PE_Array_2_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_23_io_in_psum = PE_Array_2_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_24_clock = clock;
  assign PE_Array_3_24_reset = reset;
  assign PE_Array_3_24_io_in_activate = PE_Array_3_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_24_io_in_weight = PE_Array_2_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_24_io_in_psum = PE_Array_2_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_25_clock = clock;
  assign PE_Array_3_25_reset = reset;
  assign PE_Array_3_25_io_in_activate = PE_Array_3_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_25_io_in_weight = PE_Array_2_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_25_io_in_psum = PE_Array_2_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_26_clock = clock;
  assign PE_Array_3_26_reset = reset;
  assign PE_Array_3_26_io_in_activate = PE_Array_3_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_26_io_in_weight = PE_Array_2_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_26_io_in_psum = PE_Array_2_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_27_clock = clock;
  assign PE_Array_3_27_reset = reset;
  assign PE_Array_3_27_io_in_activate = PE_Array_3_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_27_io_in_weight = PE_Array_2_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_27_io_in_psum = PE_Array_2_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_28_clock = clock;
  assign PE_Array_3_28_reset = reset;
  assign PE_Array_3_28_io_in_activate = PE_Array_3_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_28_io_in_weight = PE_Array_2_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_28_io_in_psum = PE_Array_2_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_29_clock = clock;
  assign PE_Array_3_29_reset = reset;
  assign PE_Array_3_29_io_in_activate = PE_Array_3_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_29_io_in_weight = PE_Array_2_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_29_io_in_psum = PE_Array_2_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_30_clock = clock;
  assign PE_Array_3_30_reset = reset;
  assign PE_Array_3_30_io_in_activate = PE_Array_3_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_30_io_in_weight = PE_Array_2_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_30_io_in_psum = PE_Array_2_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_31_clock = clock;
  assign PE_Array_3_31_reset = reset;
  assign PE_Array_3_31_io_in_activate = PE_Array_3_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_31_io_in_weight = PE_Array_2_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_31_io_in_psum = PE_Array_2_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_0_clock = clock;
  assign PE_Array_4_0_reset = reset;
  assign PE_Array_4_0_io_in_activate = io_activate_4; // @[DataPath.scala 11:26]
  assign PE_Array_4_0_io_in_weight = PE_Array_3_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_0_io_in_psum = PE_Array_3_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_1_clock = clock;
  assign PE_Array_4_1_reset = reset;
  assign PE_Array_4_1_io_in_activate = PE_Array_4_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_1_io_in_weight = PE_Array_3_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_1_io_in_psum = PE_Array_3_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_2_clock = clock;
  assign PE_Array_4_2_reset = reset;
  assign PE_Array_4_2_io_in_activate = PE_Array_4_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_2_io_in_weight = PE_Array_3_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_2_io_in_psum = PE_Array_3_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_3_clock = clock;
  assign PE_Array_4_3_reset = reset;
  assign PE_Array_4_3_io_in_activate = PE_Array_4_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_3_io_in_weight = PE_Array_3_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_3_io_in_psum = PE_Array_3_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_4_clock = clock;
  assign PE_Array_4_4_reset = reset;
  assign PE_Array_4_4_io_in_activate = PE_Array_4_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_4_io_in_weight = PE_Array_3_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_4_io_in_psum = PE_Array_3_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_5_clock = clock;
  assign PE_Array_4_5_reset = reset;
  assign PE_Array_4_5_io_in_activate = PE_Array_4_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_5_io_in_weight = PE_Array_3_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_5_io_in_psum = PE_Array_3_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_6_clock = clock;
  assign PE_Array_4_6_reset = reset;
  assign PE_Array_4_6_io_in_activate = PE_Array_4_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_6_io_in_weight = PE_Array_3_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_6_io_in_psum = PE_Array_3_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_7_clock = clock;
  assign PE_Array_4_7_reset = reset;
  assign PE_Array_4_7_io_in_activate = PE_Array_4_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_7_io_in_weight = PE_Array_3_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_7_io_in_psum = PE_Array_3_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_8_clock = clock;
  assign PE_Array_4_8_reset = reset;
  assign PE_Array_4_8_io_in_activate = PE_Array_4_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_8_io_in_weight = PE_Array_3_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_8_io_in_psum = PE_Array_3_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_9_clock = clock;
  assign PE_Array_4_9_reset = reset;
  assign PE_Array_4_9_io_in_activate = PE_Array_4_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_9_io_in_weight = PE_Array_3_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_9_io_in_psum = PE_Array_3_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_10_clock = clock;
  assign PE_Array_4_10_reset = reset;
  assign PE_Array_4_10_io_in_activate = PE_Array_4_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_10_io_in_weight = PE_Array_3_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_10_io_in_psum = PE_Array_3_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_11_clock = clock;
  assign PE_Array_4_11_reset = reset;
  assign PE_Array_4_11_io_in_activate = PE_Array_4_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_11_io_in_weight = PE_Array_3_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_11_io_in_psum = PE_Array_3_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_12_clock = clock;
  assign PE_Array_4_12_reset = reset;
  assign PE_Array_4_12_io_in_activate = PE_Array_4_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_12_io_in_weight = PE_Array_3_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_12_io_in_psum = PE_Array_3_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_13_clock = clock;
  assign PE_Array_4_13_reset = reset;
  assign PE_Array_4_13_io_in_activate = PE_Array_4_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_13_io_in_weight = PE_Array_3_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_13_io_in_psum = PE_Array_3_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_14_clock = clock;
  assign PE_Array_4_14_reset = reset;
  assign PE_Array_4_14_io_in_activate = PE_Array_4_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_14_io_in_weight = PE_Array_3_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_14_io_in_psum = PE_Array_3_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_15_clock = clock;
  assign PE_Array_4_15_reset = reset;
  assign PE_Array_4_15_io_in_activate = PE_Array_4_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_15_io_in_weight = PE_Array_3_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_15_io_in_psum = PE_Array_3_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_16_clock = clock;
  assign PE_Array_4_16_reset = reset;
  assign PE_Array_4_16_io_in_activate = PE_Array_4_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_16_io_in_weight = PE_Array_3_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_16_io_in_psum = PE_Array_3_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_17_clock = clock;
  assign PE_Array_4_17_reset = reset;
  assign PE_Array_4_17_io_in_activate = PE_Array_4_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_17_io_in_weight = PE_Array_3_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_17_io_in_psum = PE_Array_3_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_18_clock = clock;
  assign PE_Array_4_18_reset = reset;
  assign PE_Array_4_18_io_in_activate = PE_Array_4_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_18_io_in_weight = PE_Array_3_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_18_io_in_psum = PE_Array_3_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_19_clock = clock;
  assign PE_Array_4_19_reset = reset;
  assign PE_Array_4_19_io_in_activate = PE_Array_4_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_19_io_in_weight = PE_Array_3_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_19_io_in_psum = PE_Array_3_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_20_clock = clock;
  assign PE_Array_4_20_reset = reset;
  assign PE_Array_4_20_io_in_activate = PE_Array_4_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_20_io_in_weight = PE_Array_3_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_20_io_in_psum = PE_Array_3_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_21_clock = clock;
  assign PE_Array_4_21_reset = reset;
  assign PE_Array_4_21_io_in_activate = PE_Array_4_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_21_io_in_weight = PE_Array_3_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_21_io_in_psum = PE_Array_3_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_22_clock = clock;
  assign PE_Array_4_22_reset = reset;
  assign PE_Array_4_22_io_in_activate = PE_Array_4_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_22_io_in_weight = PE_Array_3_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_22_io_in_psum = PE_Array_3_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_23_clock = clock;
  assign PE_Array_4_23_reset = reset;
  assign PE_Array_4_23_io_in_activate = PE_Array_4_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_23_io_in_weight = PE_Array_3_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_23_io_in_psum = PE_Array_3_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_24_clock = clock;
  assign PE_Array_4_24_reset = reset;
  assign PE_Array_4_24_io_in_activate = PE_Array_4_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_24_io_in_weight = PE_Array_3_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_24_io_in_psum = PE_Array_3_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_25_clock = clock;
  assign PE_Array_4_25_reset = reset;
  assign PE_Array_4_25_io_in_activate = PE_Array_4_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_25_io_in_weight = PE_Array_3_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_25_io_in_psum = PE_Array_3_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_26_clock = clock;
  assign PE_Array_4_26_reset = reset;
  assign PE_Array_4_26_io_in_activate = PE_Array_4_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_26_io_in_weight = PE_Array_3_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_26_io_in_psum = PE_Array_3_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_27_clock = clock;
  assign PE_Array_4_27_reset = reset;
  assign PE_Array_4_27_io_in_activate = PE_Array_4_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_27_io_in_weight = PE_Array_3_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_27_io_in_psum = PE_Array_3_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_28_clock = clock;
  assign PE_Array_4_28_reset = reset;
  assign PE_Array_4_28_io_in_activate = PE_Array_4_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_28_io_in_weight = PE_Array_3_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_28_io_in_psum = PE_Array_3_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_29_clock = clock;
  assign PE_Array_4_29_reset = reset;
  assign PE_Array_4_29_io_in_activate = PE_Array_4_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_29_io_in_weight = PE_Array_3_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_29_io_in_psum = PE_Array_3_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_30_clock = clock;
  assign PE_Array_4_30_reset = reset;
  assign PE_Array_4_30_io_in_activate = PE_Array_4_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_30_io_in_weight = PE_Array_3_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_30_io_in_psum = PE_Array_3_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_31_clock = clock;
  assign PE_Array_4_31_reset = reset;
  assign PE_Array_4_31_io_in_activate = PE_Array_4_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_31_io_in_weight = PE_Array_3_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_31_io_in_psum = PE_Array_3_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_0_clock = clock;
  assign PE_Array_5_0_reset = reset;
  assign PE_Array_5_0_io_in_activate = io_activate_5; // @[DataPath.scala 11:26]
  assign PE_Array_5_0_io_in_weight = PE_Array_4_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_0_io_in_psum = PE_Array_4_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_1_clock = clock;
  assign PE_Array_5_1_reset = reset;
  assign PE_Array_5_1_io_in_activate = PE_Array_5_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_1_io_in_weight = PE_Array_4_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_1_io_in_psum = PE_Array_4_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_2_clock = clock;
  assign PE_Array_5_2_reset = reset;
  assign PE_Array_5_2_io_in_activate = PE_Array_5_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_2_io_in_weight = PE_Array_4_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_2_io_in_psum = PE_Array_4_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_3_clock = clock;
  assign PE_Array_5_3_reset = reset;
  assign PE_Array_5_3_io_in_activate = PE_Array_5_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_3_io_in_weight = PE_Array_4_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_3_io_in_psum = PE_Array_4_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_4_clock = clock;
  assign PE_Array_5_4_reset = reset;
  assign PE_Array_5_4_io_in_activate = PE_Array_5_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_4_io_in_weight = PE_Array_4_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_4_io_in_psum = PE_Array_4_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_5_clock = clock;
  assign PE_Array_5_5_reset = reset;
  assign PE_Array_5_5_io_in_activate = PE_Array_5_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_5_io_in_weight = PE_Array_4_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_5_io_in_psum = PE_Array_4_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_6_clock = clock;
  assign PE_Array_5_6_reset = reset;
  assign PE_Array_5_6_io_in_activate = PE_Array_5_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_6_io_in_weight = PE_Array_4_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_6_io_in_psum = PE_Array_4_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_7_clock = clock;
  assign PE_Array_5_7_reset = reset;
  assign PE_Array_5_7_io_in_activate = PE_Array_5_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_7_io_in_weight = PE_Array_4_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_7_io_in_psum = PE_Array_4_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_8_clock = clock;
  assign PE_Array_5_8_reset = reset;
  assign PE_Array_5_8_io_in_activate = PE_Array_5_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_8_io_in_weight = PE_Array_4_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_8_io_in_psum = PE_Array_4_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_9_clock = clock;
  assign PE_Array_5_9_reset = reset;
  assign PE_Array_5_9_io_in_activate = PE_Array_5_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_9_io_in_weight = PE_Array_4_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_9_io_in_psum = PE_Array_4_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_10_clock = clock;
  assign PE_Array_5_10_reset = reset;
  assign PE_Array_5_10_io_in_activate = PE_Array_5_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_10_io_in_weight = PE_Array_4_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_10_io_in_psum = PE_Array_4_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_11_clock = clock;
  assign PE_Array_5_11_reset = reset;
  assign PE_Array_5_11_io_in_activate = PE_Array_5_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_11_io_in_weight = PE_Array_4_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_11_io_in_psum = PE_Array_4_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_12_clock = clock;
  assign PE_Array_5_12_reset = reset;
  assign PE_Array_5_12_io_in_activate = PE_Array_5_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_12_io_in_weight = PE_Array_4_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_12_io_in_psum = PE_Array_4_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_13_clock = clock;
  assign PE_Array_5_13_reset = reset;
  assign PE_Array_5_13_io_in_activate = PE_Array_5_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_13_io_in_weight = PE_Array_4_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_13_io_in_psum = PE_Array_4_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_14_clock = clock;
  assign PE_Array_5_14_reset = reset;
  assign PE_Array_5_14_io_in_activate = PE_Array_5_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_14_io_in_weight = PE_Array_4_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_14_io_in_psum = PE_Array_4_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_15_clock = clock;
  assign PE_Array_5_15_reset = reset;
  assign PE_Array_5_15_io_in_activate = PE_Array_5_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_15_io_in_weight = PE_Array_4_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_15_io_in_psum = PE_Array_4_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_16_clock = clock;
  assign PE_Array_5_16_reset = reset;
  assign PE_Array_5_16_io_in_activate = PE_Array_5_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_16_io_in_weight = PE_Array_4_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_16_io_in_psum = PE_Array_4_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_17_clock = clock;
  assign PE_Array_5_17_reset = reset;
  assign PE_Array_5_17_io_in_activate = PE_Array_5_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_17_io_in_weight = PE_Array_4_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_17_io_in_psum = PE_Array_4_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_18_clock = clock;
  assign PE_Array_5_18_reset = reset;
  assign PE_Array_5_18_io_in_activate = PE_Array_5_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_18_io_in_weight = PE_Array_4_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_18_io_in_psum = PE_Array_4_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_19_clock = clock;
  assign PE_Array_5_19_reset = reset;
  assign PE_Array_5_19_io_in_activate = PE_Array_5_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_19_io_in_weight = PE_Array_4_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_19_io_in_psum = PE_Array_4_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_20_clock = clock;
  assign PE_Array_5_20_reset = reset;
  assign PE_Array_5_20_io_in_activate = PE_Array_5_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_20_io_in_weight = PE_Array_4_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_20_io_in_psum = PE_Array_4_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_21_clock = clock;
  assign PE_Array_5_21_reset = reset;
  assign PE_Array_5_21_io_in_activate = PE_Array_5_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_21_io_in_weight = PE_Array_4_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_21_io_in_psum = PE_Array_4_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_22_clock = clock;
  assign PE_Array_5_22_reset = reset;
  assign PE_Array_5_22_io_in_activate = PE_Array_5_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_22_io_in_weight = PE_Array_4_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_22_io_in_psum = PE_Array_4_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_23_clock = clock;
  assign PE_Array_5_23_reset = reset;
  assign PE_Array_5_23_io_in_activate = PE_Array_5_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_23_io_in_weight = PE_Array_4_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_23_io_in_psum = PE_Array_4_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_24_clock = clock;
  assign PE_Array_5_24_reset = reset;
  assign PE_Array_5_24_io_in_activate = PE_Array_5_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_24_io_in_weight = PE_Array_4_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_24_io_in_psum = PE_Array_4_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_25_clock = clock;
  assign PE_Array_5_25_reset = reset;
  assign PE_Array_5_25_io_in_activate = PE_Array_5_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_25_io_in_weight = PE_Array_4_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_25_io_in_psum = PE_Array_4_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_26_clock = clock;
  assign PE_Array_5_26_reset = reset;
  assign PE_Array_5_26_io_in_activate = PE_Array_5_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_26_io_in_weight = PE_Array_4_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_26_io_in_psum = PE_Array_4_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_27_clock = clock;
  assign PE_Array_5_27_reset = reset;
  assign PE_Array_5_27_io_in_activate = PE_Array_5_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_27_io_in_weight = PE_Array_4_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_27_io_in_psum = PE_Array_4_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_28_clock = clock;
  assign PE_Array_5_28_reset = reset;
  assign PE_Array_5_28_io_in_activate = PE_Array_5_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_28_io_in_weight = PE_Array_4_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_28_io_in_psum = PE_Array_4_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_29_clock = clock;
  assign PE_Array_5_29_reset = reset;
  assign PE_Array_5_29_io_in_activate = PE_Array_5_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_29_io_in_weight = PE_Array_4_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_29_io_in_psum = PE_Array_4_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_30_clock = clock;
  assign PE_Array_5_30_reset = reset;
  assign PE_Array_5_30_io_in_activate = PE_Array_5_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_30_io_in_weight = PE_Array_4_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_30_io_in_psum = PE_Array_4_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_31_clock = clock;
  assign PE_Array_5_31_reset = reset;
  assign PE_Array_5_31_io_in_activate = PE_Array_5_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_31_io_in_weight = PE_Array_4_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_31_io_in_psum = PE_Array_4_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_0_clock = clock;
  assign PE_Array_6_0_reset = reset;
  assign PE_Array_6_0_io_in_activate = io_activate_6; // @[DataPath.scala 11:26]
  assign PE_Array_6_0_io_in_weight = PE_Array_5_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_0_io_in_psum = PE_Array_5_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_1_clock = clock;
  assign PE_Array_6_1_reset = reset;
  assign PE_Array_6_1_io_in_activate = PE_Array_6_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_1_io_in_weight = PE_Array_5_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_1_io_in_psum = PE_Array_5_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_2_clock = clock;
  assign PE_Array_6_2_reset = reset;
  assign PE_Array_6_2_io_in_activate = PE_Array_6_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_2_io_in_weight = PE_Array_5_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_2_io_in_psum = PE_Array_5_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_3_clock = clock;
  assign PE_Array_6_3_reset = reset;
  assign PE_Array_6_3_io_in_activate = PE_Array_6_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_3_io_in_weight = PE_Array_5_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_3_io_in_psum = PE_Array_5_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_4_clock = clock;
  assign PE_Array_6_4_reset = reset;
  assign PE_Array_6_4_io_in_activate = PE_Array_6_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_4_io_in_weight = PE_Array_5_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_4_io_in_psum = PE_Array_5_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_5_clock = clock;
  assign PE_Array_6_5_reset = reset;
  assign PE_Array_6_5_io_in_activate = PE_Array_6_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_5_io_in_weight = PE_Array_5_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_5_io_in_psum = PE_Array_5_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_6_clock = clock;
  assign PE_Array_6_6_reset = reset;
  assign PE_Array_6_6_io_in_activate = PE_Array_6_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_6_io_in_weight = PE_Array_5_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_6_io_in_psum = PE_Array_5_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_7_clock = clock;
  assign PE_Array_6_7_reset = reset;
  assign PE_Array_6_7_io_in_activate = PE_Array_6_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_7_io_in_weight = PE_Array_5_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_7_io_in_psum = PE_Array_5_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_8_clock = clock;
  assign PE_Array_6_8_reset = reset;
  assign PE_Array_6_8_io_in_activate = PE_Array_6_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_8_io_in_weight = PE_Array_5_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_8_io_in_psum = PE_Array_5_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_9_clock = clock;
  assign PE_Array_6_9_reset = reset;
  assign PE_Array_6_9_io_in_activate = PE_Array_6_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_9_io_in_weight = PE_Array_5_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_9_io_in_psum = PE_Array_5_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_10_clock = clock;
  assign PE_Array_6_10_reset = reset;
  assign PE_Array_6_10_io_in_activate = PE_Array_6_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_10_io_in_weight = PE_Array_5_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_10_io_in_psum = PE_Array_5_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_11_clock = clock;
  assign PE_Array_6_11_reset = reset;
  assign PE_Array_6_11_io_in_activate = PE_Array_6_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_11_io_in_weight = PE_Array_5_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_11_io_in_psum = PE_Array_5_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_12_clock = clock;
  assign PE_Array_6_12_reset = reset;
  assign PE_Array_6_12_io_in_activate = PE_Array_6_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_12_io_in_weight = PE_Array_5_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_12_io_in_psum = PE_Array_5_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_13_clock = clock;
  assign PE_Array_6_13_reset = reset;
  assign PE_Array_6_13_io_in_activate = PE_Array_6_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_13_io_in_weight = PE_Array_5_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_13_io_in_psum = PE_Array_5_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_14_clock = clock;
  assign PE_Array_6_14_reset = reset;
  assign PE_Array_6_14_io_in_activate = PE_Array_6_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_14_io_in_weight = PE_Array_5_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_14_io_in_psum = PE_Array_5_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_15_clock = clock;
  assign PE_Array_6_15_reset = reset;
  assign PE_Array_6_15_io_in_activate = PE_Array_6_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_15_io_in_weight = PE_Array_5_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_15_io_in_psum = PE_Array_5_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_16_clock = clock;
  assign PE_Array_6_16_reset = reset;
  assign PE_Array_6_16_io_in_activate = PE_Array_6_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_16_io_in_weight = PE_Array_5_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_16_io_in_psum = PE_Array_5_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_17_clock = clock;
  assign PE_Array_6_17_reset = reset;
  assign PE_Array_6_17_io_in_activate = PE_Array_6_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_17_io_in_weight = PE_Array_5_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_17_io_in_psum = PE_Array_5_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_18_clock = clock;
  assign PE_Array_6_18_reset = reset;
  assign PE_Array_6_18_io_in_activate = PE_Array_6_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_18_io_in_weight = PE_Array_5_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_18_io_in_psum = PE_Array_5_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_19_clock = clock;
  assign PE_Array_6_19_reset = reset;
  assign PE_Array_6_19_io_in_activate = PE_Array_6_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_19_io_in_weight = PE_Array_5_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_19_io_in_psum = PE_Array_5_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_20_clock = clock;
  assign PE_Array_6_20_reset = reset;
  assign PE_Array_6_20_io_in_activate = PE_Array_6_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_20_io_in_weight = PE_Array_5_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_20_io_in_psum = PE_Array_5_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_21_clock = clock;
  assign PE_Array_6_21_reset = reset;
  assign PE_Array_6_21_io_in_activate = PE_Array_6_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_21_io_in_weight = PE_Array_5_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_21_io_in_psum = PE_Array_5_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_22_clock = clock;
  assign PE_Array_6_22_reset = reset;
  assign PE_Array_6_22_io_in_activate = PE_Array_6_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_22_io_in_weight = PE_Array_5_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_22_io_in_psum = PE_Array_5_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_23_clock = clock;
  assign PE_Array_6_23_reset = reset;
  assign PE_Array_6_23_io_in_activate = PE_Array_6_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_23_io_in_weight = PE_Array_5_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_23_io_in_psum = PE_Array_5_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_24_clock = clock;
  assign PE_Array_6_24_reset = reset;
  assign PE_Array_6_24_io_in_activate = PE_Array_6_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_24_io_in_weight = PE_Array_5_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_24_io_in_psum = PE_Array_5_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_25_clock = clock;
  assign PE_Array_6_25_reset = reset;
  assign PE_Array_6_25_io_in_activate = PE_Array_6_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_25_io_in_weight = PE_Array_5_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_25_io_in_psum = PE_Array_5_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_26_clock = clock;
  assign PE_Array_6_26_reset = reset;
  assign PE_Array_6_26_io_in_activate = PE_Array_6_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_26_io_in_weight = PE_Array_5_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_26_io_in_psum = PE_Array_5_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_27_clock = clock;
  assign PE_Array_6_27_reset = reset;
  assign PE_Array_6_27_io_in_activate = PE_Array_6_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_27_io_in_weight = PE_Array_5_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_27_io_in_psum = PE_Array_5_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_28_clock = clock;
  assign PE_Array_6_28_reset = reset;
  assign PE_Array_6_28_io_in_activate = PE_Array_6_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_28_io_in_weight = PE_Array_5_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_28_io_in_psum = PE_Array_5_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_29_clock = clock;
  assign PE_Array_6_29_reset = reset;
  assign PE_Array_6_29_io_in_activate = PE_Array_6_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_29_io_in_weight = PE_Array_5_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_29_io_in_psum = PE_Array_5_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_30_clock = clock;
  assign PE_Array_6_30_reset = reset;
  assign PE_Array_6_30_io_in_activate = PE_Array_6_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_30_io_in_weight = PE_Array_5_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_30_io_in_psum = PE_Array_5_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_31_clock = clock;
  assign PE_Array_6_31_reset = reset;
  assign PE_Array_6_31_io_in_activate = PE_Array_6_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_31_io_in_weight = PE_Array_5_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_31_io_in_psum = PE_Array_5_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_0_clock = clock;
  assign PE_Array_7_0_reset = reset;
  assign PE_Array_7_0_io_in_activate = io_activate_7; // @[DataPath.scala 11:26]
  assign PE_Array_7_0_io_in_weight = PE_Array_6_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_0_io_in_psum = PE_Array_6_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_1_clock = clock;
  assign PE_Array_7_1_reset = reset;
  assign PE_Array_7_1_io_in_activate = PE_Array_7_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_1_io_in_weight = PE_Array_6_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_1_io_in_psum = PE_Array_6_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_2_clock = clock;
  assign PE_Array_7_2_reset = reset;
  assign PE_Array_7_2_io_in_activate = PE_Array_7_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_2_io_in_weight = PE_Array_6_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_2_io_in_psum = PE_Array_6_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_3_clock = clock;
  assign PE_Array_7_3_reset = reset;
  assign PE_Array_7_3_io_in_activate = PE_Array_7_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_3_io_in_weight = PE_Array_6_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_3_io_in_psum = PE_Array_6_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_4_clock = clock;
  assign PE_Array_7_4_reset = reset;
  assign PE_Array_7_4_io_in_activate = PE_Array_7_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_4_io_in_weight = PE_Array_6_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_4_io_in_psum = PE_Array_6_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_5_clock = clock;
  assign PE_Array_7_5_reset = reset;
  assign PE_Array_7_5_io_in_activate = PE_Array_7_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_5_io_in_weight = PE_Array_6_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_5_io_in_psum = PE_Array_6_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_6_clock = clock;
  assign PE_Array_7_6_reset = reset;
  assign PE_Array_7_6_io_in_activate = PE_Array_7_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_6_io_in_weight = PE_Array_6_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_6_io_in_psum = PE_Array_6_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_7_clock = clock;
  assign PE_Array_7_7_reset = reset;
  assign PE_Array_7_7_io_in_activate = PE_Array_7_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_7_io_in_weight = PE_Array_6_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_7_io_in_psum = PE_Array_6_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_8_clock = clock;
  assign PE_Array_7_8_reset = reset;
  assign PE_Array_7_8_io_in_activate = PE_Array_7_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_8_io_in_weight = PE_Array_6_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_8_io_in_psum = PE_Array_6_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_9_clock = clock;
  assign PE_Array_7_9_reset = reset;
  assign PE_Array_7_9_io_in_activate = PE_Array_7_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_9_io_in_weight = PE_Array_6_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_9_io_in_psum = PE_Array_6_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_10_clock = clock;
  assign PE_Array_7_10_reset = reset;
  assign PE_Array_7_10_io_in_activate = PE_Array_7_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_10_io_in_weight = PE_Array_6_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_10_io_in_psum = PE_Array_6_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_11_clock = clock;
  assign PE_Array_7_11_reset = reset;
  assign PE_Array_7_11_io_in_activate = PE_Array_7_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_11_io_in_weight = PE_Array_6_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_11_io_in_psum = PE_Array_6_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_12_clock = clock;
  assign PE_Array_7_12_reset = reset;
  assign PE_Array_7_12_io_in_activate = PE_Array_7_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_12_io_in_weight = PE_Array_6_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_12_io_in_psum = PE_Array_6_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_13_clock = clock;
  assign PE_Array_7_13_reset = reset;
  assign PE_Array_7_13_io_in_activate = PE_Array_7_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_13_io_in_weight = PE_Array_6_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_13_io_in_psum = PE_Array_6_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_14_clock = clock;
  assign PE_Array_7_14_reset = reset;
  assign PE_Array_7_14_io_in_activate = PE_Array_7_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_14_io_in_weight = PE_Array_6_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_14_io_in_psum = PE_Array_6_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_15_clock = clock;
  assign PE_Array_7_15_reset = reset;
  assign PE_Array_7_15_io_in_activate = PE_Array_7_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_15_io_in_weight = PE_Array_6_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_15_io_in_psum = PE_Array_6_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_16_clock = clock;
  assign PE_Array_7_16_reset = reset;
  assign PE_Array_7_16_io_in_activate = PE_Array_7_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_16_io_in_weight = PE_Array_6_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_16_io_in_psum = PE_Array_6_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_17_clock = clock;
  assign PE_Array_7_17_reset = reset;
  assign PE_Array_7_17_io_in_activate = PE_Array_7_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_17_io_in_weight = PE_Array_6_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_17_io_in_psum = PE_Array_6_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_18_clock = clock;
  assign PE_Array_7_18_reset = reset;
  assign PE_Array_7_18_io_in_activate = PE_Array_7_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_18_io_in_weight = PE_Array_6_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_18_io_in_psum = PE_Array_6_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_19_clock = clock;
  assign PE_Array_7_19_reset = reset;
  assign PE_Array_7_19_io_in_activate = PE_Array_7_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_19_io_in_weight = PE_Array_6_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_19_io_in_psum = PE_Array_6_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_20_clock = clock;
  assign PE_Array_7_20_reset = reset;
  assign PE_Array_7_20_io_in_activate = PE_Array_7_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_20_io_in_weight = PE_Array_6_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_20_io_in_psum = PE_Array_6_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_21_clock = clock;
  assign PE_Array_7_21_reset = reset;
  assign PE_Array_7_21_io_in_activate = PE_Array_7_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_21_io_in_weight = PE_Array_6_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_21_io_in_psum = PE_Array_6_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_22_clock = clock;
  assign PE_Array_7_22_reset = reset;
  assign PE_Array_7_22_io_in_activate = PE_Array_7_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_22_io_in_weight = PE_Array_6_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_22_io_in_psum = PE_Array_6_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_23_clock = clock;
  assign PE_Array_7_23_reset = reset;
  assign PE_Array_7_23_io_in_activate = PE_Array_7_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_23_io_in_weight = PE_Array_6_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_23_io_in_psum = PE_Array_6_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_24_clock = clock;
  assign PE_Array_7_24_reset = reset;
  assign PE_Array_7_24_io_in_activate = PE_Array_7_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_24_io_in_weight = PE_Array_6_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_24_io_in_psum = PE_Array_6_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_25_clock = clock;
  assign PE_Array_7_25_reset = reset;
  assign PE_Array_7_25_io_in_activate = PE_Array_7_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_25_io_in_weight = PE_Array_6_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_25_io_in_psum = PE_Array_6_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_26_clock = clock;
  assign PE_Array_7_26_reset = reset;
  assign PE_Array_7_26_io_in_activate = PE_Array_7_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_26_io_in_weight = PE_Array_6_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_26_io_in_psum = PE_Array_6_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_27_clock = clock;
  assign PE_Array_7_27_reset = reset;
  assign PE_Array_7_27_io_in_activate = PE_Array_7_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_27_io_in_weight = PE_Array_6_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_27_io_in_psum = PE_Array_6_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_28_clock = clock;
  assign PE_Array_7_28_reset = reset;
  assign PE_Array_7_28_io_in_activate = PE_Array_7_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_28_io_in_weight = PE_Array_6_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_28_io_in_psum = PE_Array_6_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_29_clock = clock;
  assign PE_Array_7_29_reset = reset;
  assign PE_Array_7_29_io_in_activate = PE_Array_7_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_29_io_in_weight = PE_Array_6_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_29_io_in_psum = PE_Array_6_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_30_clock = clock;
  assign PE_Array_7_30_reset = reset;
  assign PE_Array_7_30_io_in_activate = PE_Array_7_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_30_io_in_weight = PE_Array_6_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_30_io_in_psum = PE_Array_6_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_31_clock = clock;
  assign PE_Array_7_31_reset = reset;
  assign PE_Array_7_31_io_in_activate = PE_Array_7_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_31_io_in_weight = PE_Array_6_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_31_io_in_psum = PE_Array_6_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_0_clock = clock;
  assign PE_Array_8_0_reset = reset;
  assign PE_Array_8_0_io_in_activate = io_activate_8; // @[DataPath.scala 11:26]
  assign PE_Array_8_0_io_in_weight = PE_Array_7_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_0_io_in_psum = PE_Array_7_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_1_clock = clock;
  assign PE_Array_8_1_reset = reset;
  assign PE_Array_8_1_io_in_activate = PE_Array_8_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_1_io_in_weight = PE_Array_7_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_1_io_in_psum = PE_Array_7_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_2_clock = clock;
  assign PE_Array_8_2_reset = reset;
  assign PE_Array_8_2_io_in_activate = PE_Array_8_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_2_io_in_weight = PE_Array_7_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_2_io_in_psum = PE_Array_7_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_3_clock = clock;
  assign PE_Array_8_3_reset = reset;
  assign PE_Array_8_3_io_in_activate = PE_Array_8_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_3_io_in_weight = PE_Array_7_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_3_io_in_psum = PE_Array_7_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_4_clock = clock;
  assign PE_Array_8_4_reset = reset;
  assign PE_Array_8_4_io_in_activate = PE_Array_8_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_4_io_in_weight = PE_Array_7_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_4_io_in_psum = PE_Array_7_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_5_clock = clock;
  assign PE_Array_8_5_reset = reset;
  assign PE_Array_8_5_io_in_activate = PE_Array_8_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_5_io_in_weight = PE_Array_7_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_5_io_in_psum = PE_Array_7_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_6_clock = clock;
  assign PE_Array_8_6_reset = reset;
  assign PE_Array_8_6_io_in_activate = PE_Array_8_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_6_io_in_weight = PE_Array_7_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_6_io_in_psum = PE_Array_7_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_7_clock = clock;
  assign PE_Array_8_7_reset = reset;
  assign PE_Array_8_7_io_in_activate = PE_Array_8_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_7_io_in_weight = PE_Array_7_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_7_io_in_psum = PE_Array_7_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_8_clock = clock;
  assign PE_Array_8_8_reset = reset;
  assign PE_Array_8_8_io_in_activate = PE_Array_8_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_8_io_in_weight = PE_Array_7_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_8_io_in_psum = PE_Array_7_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_9_clock = clock;
  assign PE_Array_8_9_reset = reset;
  assign PE_Array_8_9_io_in_activate = PE_Array_8_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_9_io_in_weight = PE_Array_7_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_9_io_in_psum = PE_Array_7_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_10_clock = clock;
  assign PE_Array_8_10_reset = reset;
  assign PE_Array_8_10_io_in_activate = PE_Array_8_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_10_io_in_weight = PE_Array_7_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_10_io_in_psum = PE_Array_7_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_11_clock = clock;
  assign PE_Array_8_11_reset = reset;
  assign PE_Array_8_11_io_in_activate = PE_Array_8_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_11_io_in_weight = PE_Array_7_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_11_io_in_psum = PE_Array_7_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_12_clock = clock;
  assign PE_Array_8_12_reset = reset;
  assign PE_Array_8_12_io_in_activate = PE_Array_8_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_12_io_in_weight = PE_Array_7_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_12_io_in_psum = PE_Array_7_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_13_clock = clock;
  assign PE_Array_8_13_reset = reset;
  assign PE_Array_8_13_io_in_activate = PE_Array_8_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_13_io_in_weight = PE_Array_7_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_13_io_in_psum = PE_Array_7_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_14_clock = clock;
  assign PE_Array_8_14_reset = reset;
  assign PE_Array_8_14_io_in_activate = PE_Array_8_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_14_io_in_weight = PE_Array_7_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_14_io_in_psum = PE_Array_7_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_15_clock = clock;
  assign PE_Array_8_15_reset = reset;
  assign PE_Array_8_15_io_in_activate = PE_Array_8_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_15_io_in_weight = PE_Array_7_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_15_io_in_psum = PE_Array_7_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_16_clock = clock;
  assign PE_Array_8_16_reset = reset;
  assign PE_Array_8_16_io_in_activate = PE_Array_8_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_16_io_in_weight = PE_Array_7_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_16_io_in_psum = PE_Array_7_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_17_clock = clock;
  assign PE_Array_8_17_reset = reset;
  assign PE_Array_8_17_io_in_activate = PE_Array_8_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_17_io_in_weight = PE_Array_7_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_17_io_in_psum = PE_Array_7_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_18_clock = clock;
  assign PE_Array_8_18_reset = reset;
  assign PE_Array_8_18_io_in_activate = PE_Array_8_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_18_io_in_weight = PE_Array_7_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_18_io_in_psum = PE_Array_7_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_19_clock = clock;
  assign PE_Array_8_19_reset = reset;
  assign PE_Array_8_19_io_in_activate = PE_Array_8_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_19_io_in_weight = PE_Array_7_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_19_io_in_psum = PE_Array_7_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_20_clock = clock;
  assign PE_Array_8_20_reset = reset;
  assign PE_Array_8_20_io_in_activate = PE_Array_8_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_20_io_in_weight = PE_Array_7_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_20_io_in_psum = PE_Array_7_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_21_clock = clock;
  assign PE_Array_8_21_reset = reset;
  assign PE_Array_8_21_io_in_activate = PE_Array_8_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_21_io_in_weight = PE_Array_7_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_21_io_in_psum = PE_Array_7_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_22_clock = clock;
  assign PE_Array_8_22_reset = reset;
  assign PE_Array_8_22_io_in_activate = PE_Array_8_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_22_io_in_weight = PE_Array_7_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_22_io_in_psum = PE_Array_7_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_23_clock = clock;
  assign PE_Array_8_23_reset = reset;
  assign PE_Array_8_23_io_in_activate = PE_Array_8_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_23_io_in_weight = PE_Array_7_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_23_io_in_psum = PE_Array_7_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_24_clock = clock;
  assign PE_Array_8_24_reset = reset;
  assign PE_Array_8_24_io_in_activate = PE_Array_8_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_24_io_in_weight = PE_Array_7_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_24_io_in_psum = PE_Array_7_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_25_clock = clock;
  assign PE_Array_8_25_reset = reset;
  assign PE_Array_8_25_io_in_activate = PE_Array_8_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_25_io_in_weight = PE_Array_7_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_25_io_in_psum = PE_Array_7_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_26_clock = clock;
  assign PE_Array_8_26_reset = reset;
  assign PE_Array_8_26_io_in_activate = PE_Array_8_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_26_io_in_weight = PE_Array_7_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_26_io_in_psum = PE_Array_7_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_27_clock = clock;
  assign PE_Array_8_27_reset = reset;
  assign PE_Array_8_27_io_in_activate = PE_Array_8_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_27_io_in_weight = PE_Array_7_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_27_io_in_psum = PE_Array_7_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_28_clock = clock;
  assign PE_Array_8_28_reset = reset;
  assign PE_Array_8_28_io_in_activate = PE_Array_8_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_28_io_in_weight = PE_Array_7_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_28_io_in_psum = PE_Array_7_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_29_clock = clock;
  assign PE_Array_8_29_reset = reset;
  assign PE_Array_8_29_io_in_activate = PE_Array_8_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_29_io_in_weight = PE_Array_7_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_29_io_in_psum = PE_Array_7_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_30_clock = clock;
  assign PE_Array_8_30_reset = reset;
  assign PE_Array_8_30_io_in_activate = PE_Array_8_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_30_io_in_weight = PE_Array_7_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_30_io_in_psum = PE_Array_7_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_8_31_clock = clock;
  assign PE_Array_8_31_reset = reset;
  assign PE_Array_8_31_io_in_activate = PE_Array_8_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_8_31_io_in_weight = PE_Array_7_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_8_31_io_in_psum = PE_Array_7_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_8_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_8_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_0_clock = clock;
  assign PE_Array_9_0_reset = reset;
  assign PE_Array_9_0_io_in_activate = io_activate_9; // @[DataPath.scala 11:26]
  assign PE_Array_9_0_io_in_weight = PE_Array_8_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_0_io_in_psum = PE_Array_8_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_1_clock = clock;
  assign PE_Array_9_1_reset = reset;
  assign PE_Array_9_1_io_in_activate = PE_Array_9_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_1_io_in_weight = PE_Array_8_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_1_io_in_psum = PE_Array_8_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_2_clock = clock;
  assign PE_Array_9_2_reset = reset;
  assign PE_Array_9_2_io_in_activate = PE_Array_9_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_2_io_in_weight = PE_Array_8_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_2_io_in_psum = PE_Array_8_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_3_clock = clock;
  assign PE_Array_9_3_reset = reset;
  assign PE_Array_9_3_io_in_activate = PE_Array_9_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_3_io_in_weight = PE_Array_8_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_3_io_in_psum = PE_Array_8_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_4_clock = clock;
  assign PE_Array_9_4_reset = reset;
  assign PE_Array_9_4_io_in_activate = PE_Array_9_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_4_io_in_weight = PE_Array_8_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_4_io_in_psum = PE_Array_8_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_5_clock = clock;
  assign PE_Array_9_5_reset = reset;
  assign PE_Array_9_5_io_in_activate = PE_Array_9_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_5_io_in_weight = PE_Array_8_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_5_io_in_psum = PE_Array_8_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_6_clock = clock;
  assign PE_Array_9_6_reset = reset;
  assign PE_Array_9_6_io_in_activate = PE_Array_9_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_6_io_in_weight = PE_Array_8_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_6_io_in_psum = PE_Array_8_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_7_clock = clock;
  assign PE_Array_9_7_reset = reset;
  assign PE_Array_9_7_io_in_activate = PE_Array_9_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_7_io_in_weight = PE_Array_8_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_7_io_in_psum = PE_Array_8_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_8_clock = clock;
  assign PE_Array_9_8_reset = reset;
  assign PE_Array_9_8_io_in_activate = PE_Array_9_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_8_io_in_weight = PE_Array_8_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_8_io_in_psum = PE_Array_8_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_9_clock = clock;
  assign PE_Array_9_9_reset = reset;
  assign PE_Array_9_9_io_in_activate = PE_Array_9_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_9_io_in_weight = PE_Array_8_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_9_io_in_psum = PE_Array_8_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_10_clock = clock;
  assign PE_Array_9_10_reset = reset;
  assign PE_Array_9_10_io_in_activate = PE_Array_9_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_10_io_in_weight = PE_Array_8_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_10_io_in_psum = PE_Array_8_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_11_clock = clock;
  assign PE_Array_9_11_reset = reset;
  assign PE_Array_9_11_io_in_activate = PE_Array_9_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_11_io_in_weight = PE_Array_8_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_11_io_in_psum = PE_Array_8_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_12_clock = clock;
  assign PE_Array_9_12_reset = reset;
  assign PE_Array_9_12_io_in_activate = PE_Array_9_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_12_io_in_weight = PE_Array_8_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_12_io_in_psum = PE_Array_8_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_13_clock = clock;
  assign PE_Array_9_13_reset = reset;
  assign PE_Array_9_13_io_in_activate = PE_Array_9_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_13_io_in_weight = PE_Array_8_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_13_io_in_psum = PE_Array_8_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_14_clock = clock;
  assign PE_Array_9_14_reset = reset;
  assign PE_Array_9_14_io_in_activate = PE_Array_9_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_14_io_in_weight = PE_Array_8_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_14_io_in_psum = PE_Array_8_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_15_clock = clock;
  assign PE_Array_9_15_reset = reset;
  assign PE_Array_9_15_io_in_activate = PE_Array_9_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_15_io_in_weight = PE_Array_8_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_15_io_in_psum = PE_Array_8_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_16_clock = clock;
  assign PE_Array_9_16_reset = reset;
  assign PE_Array_9_16_io_in_activate = PE_Array_9_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_16_io_in_weight = PE_Array_8_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_16_io_in_psum = PE_Array_8_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_17_clock = clock;
  assign PE_Array_9_17_reset = reset;
  assign PE_Array_9_17_io_in_activate = PE_Array_9_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_17_io_in_weight = PE_Array_8_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_17_io_in_psum = PE_Array_8_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_18_clock = clock;
  assign PE_Array_9_18_reset = reset;
  assign PE_Array_9_18_io_in_activate = PE_Array_9_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_18_io_in_weight = PE_Array_8_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_18_io_in_psum = PE_Array_8_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_19_clock = clock;
  assign PE_Array_9_19_reset = reset;
  assign PE_Array_9_19_io_in_activate = PE_Array_9_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_19_io_in_weight = PE_Array_8_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_19_io_in_psum = PE_Array_8_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_20_clock = clock;
  assign PE_Array_9_20_reset = reset;
  assign PE_Array_9_20_io_in_activate = PE_Array_9_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_20_io_in_weight = PE_Array_8_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_20_io_in_psum = PE_Array_8_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_21_clock = clock;
  assign PE_Array_9_21_reset = reset;
  assign PE_Array_9_21_io_in_activate = PE_Array_9_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_21_io_in_weight = PE_Array_8_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_21_io_in_psum = PE_Array_8_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_22_clock = clock;
  assign PE_Array_9_22_reset = reset;
  assign PE_Array_9_22_io_in_activate = PE_Array_9_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_22_io_in_weight = PE_Array_8_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_22_io_in_psum = PE_Array_8_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_23_clock = clock;
  assign PE_Array_9_23_reset = reset;
  assign PE_Array_9_23_io_in_activate = PE_Array_9_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_23_io_in_weight = PE_Array_8_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_23_io_in_psum = PE_Array_8_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_24_clock = clock;
  assign PE_Array_9_24_reset = reset;
  assign PE_Array_9_24_io_in_activate = PE_Array_9_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_24_io_in_weight = PE_Array_8_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_24_io_in_psum = PE_Array_8_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_25_clock = clock;
  assign PE_Array_9_25_reset = reset;
  assign PE_Array_9_25_io_in_activate = PE_Array_9_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_25_io_in_weight = PE_Array_8_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_25_io_in_psum = PE_Array_8_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_26_clock = clock;
  assign PE_Array_9_26_reset = reset;
  assign PE_Array_9_26_io_in_activate = PE_Array_9_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_26_io_in_weight = PE_Array_8_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_26_io_in_psum = PE_Array_8_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_27_clock = clock;
  assign PE_Array_9_27_reset = reset;
  assign PE_Array_9_27_io_in_activate = PE_Array_9_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_27_io_in_weight = PE_Array_8_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_27_io_in_psum = PE_Array_8_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_28_clock = clock;
  assign PE_Array_9_28_reset = reset;
  assign PE_Array_9_28_io_in_activate = PE_Array_9_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_28_io_in_weight = PE_Array_8_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_28_io_in_psum = PE_Array_8_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_29_clock = clock;
  assign PE_Array_9_29_reset = reset;
  assign PE_Array_9_29_io_in_activate = PE_Array_9_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_29_io_in_weight = PE_Array_8_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_29_io_in_psum = PE_Array_8_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_30_clock = clock;
  assign PE_Array_9_30_reset = reset;
  assign PE_Array_9_30_io_in_activate = PE_Array_9_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_30_io_in_weight = PE_Array_8_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_30_io_in_psum = PE_Array_8_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_9_31_clock = clock;
  assign PE_Array_9_31_reset = reset;
  assign PE_Array_9_31_io_in_activate = PE_Array_9_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_9_31_io_in_weight = PE_Array_8_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_9_31_io_in_psum = PE_Array_8_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_9_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_9_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_0_clock = clock;
  assign PE_Array_10_0_reset = reset;
  assign PE_Array_10_0_io_in_activate = io_activate_10; // @[DataPath.scala 11:26]
  assign PE_Array_10_0_io_in_weight = PE_Array_9_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_0_io_in_psum = PE_Array_9_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_1_clock = clock;
  assign PE_Array_10_1_reset = reset;
  assign PE_Array_10_1_io_in_activate = PE_Array_10_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_1_io_in_weight = PE_Array_9_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_1_io_in_psum = PE_Array_9_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_2_clock = clock;
  assign PE_Array_10_2_reset = reset;
  assign PE_Array_10_2_io_in_activate = PE_Array_10_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_2_io_in_weight = PE_Array_9_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_2_io_in_psum = PE_Array_9_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_3_clock = clock;
  assign PE_Array_10_3_reset = reset;
  assign PE_Array_10_3_io_in_activate = PE_Array_10_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_3_io_in_weight = PE_Array_9_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_3_io_in_psum = PE_Array_9_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_4_clock = clock;
  assign PE_Array_10_4_reset = reset;
  assign PE_Array_10_4_io_in_activate = PE_Array_10_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_4_io_in_weight = PE_Array_9_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_4_io_in_psum = PE_Array_9_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_5_clock = clock;
  assign PE_Array_10_5_reset = reset;
  assign PE_Array_10_5_io_in_activate = PE_Array_10_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_5_io_in_weight = PE_Array_9_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_5_io_in_psum = PE_Array_9_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_6_clock = clock;
  assign PE_Array_10_6_reset = reset;
  assign PE_Array_10_6_io_in_activate = PE_Array_10_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_6_io_in_weight = PE_Array_9_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_6_io_in_psum = PE_Array_9_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_7_clock = clock;
  assign PE_Array_10_7_reset = reset;
  assign PE_Array_10_7_io_in_activate = PE_Array_10_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_7_io_in_weight = PE_Array_9_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_7_io_in_psum = PE_Array_9_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_8_clock = clock;
  assign PE_Array_10_8_reset = reset;
  assign PE_Array_10_8_io_in_activate = PE_Array_10_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_8_io_in_weight = PE_Array_9_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_8_io_in_psum = PE_Array_9_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_9_clock = clock;
  assign PE_Array_10_9_reset = reset;
  assign PE_Array_10_9_io_in_activate = PE_Array_10_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_9_io_in_weight = PE_Array_9_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_9_io_in_psum = PE_Array_9_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_10_clock = clock;
  assign PE_Array_10_10_reset = reset;
  assign PE_Array_10_10_io_in_activate = PE_Array_10_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_10_io_in_weight = PE_Array_9_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_10_io_in_psum = PE_Array_9_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_11_clock = clock;
  assign PE_Array_10_11_reset = reset;
  assign PE_Array_10_11_io_in_activate = PE_Array_10_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_11_io_in_weight = PE_Array_9_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_11_io_in_psum = PE_Array_9_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_12_clock = clock;
  assign PE_Array_10_12_reset = reset;
  assign PE_Array_10_12_io_in_activate = PE_Array_10_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_12_io_in_weight = PE_Array_9_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_12_io_in_psum = PE_Array_9_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_13_clock = clock;
  assign PE_Array_10_13_reset = reset;
  assign PE_Array_10_13_io_in_activate = PE_Array_10_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_13_io_in_weight = PE_Array_9_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_13_io_in_psum = PE_Array_9_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_14_clock = clock;
  assign PE_Array_10_14_reset = reset;
  assign PE_Array_10_14_io_in_activate = PE_Array_10_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_14_io_in_weight = PE_Array_9_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_14_io_in_psum = PE_Array_9_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_15_clock = clock;
  assign PE_Array_10_15_reset = reset;
  assign PE_Array_10_15_io_in_activate = PE_Array_10_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_15_io_in_weight = PE_Array_9_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_15_io_in_psum = PE_Array_9_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_16_clock = clock;
  assign PE_Array_10_16_reset = reset;
  assign PE_Array_10_16_io_in_activate = PE_Array_10_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_16_io_in_weight = PE_Array_9_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_16_io_in_psum = PE_Array_9_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_17_clock = clock;
  assign PE_Array_10_17_reset = reset;
  assign PE_Array_10_17_io_in_activate = PE_Array_10_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_17_io_in_weight = PE_Array_9_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_17_io_in_psum = PE_Array_9_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_18_clock = clock;
  assign PE_Array_10_18_reset = reset;
  assign PE_Array_10_18_io_in_activate = PE_Array_10_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_18_io_in_weight = PE_Array_9_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_18_io_in_psum = PE_Array_9_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_19_clock = clock;
  assign PE_Array_10_19_reset = reset;
  assign PE_Array_10_19_io_in_activate = PE_Array_10_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_19_io_in_weight = PE_Array_9_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_19_io_in_psum = PE_Array_9_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_20_clock = clock;
  assign PE_Array_10_20_reset = reset;
  assign PE_Array_10_20_io_in_activate = PE_Array_10_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_20_io_in_weight = PE_Array_9_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_20_io_in_psum = PE_Array_9_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_21_clock = clock;
  assign PE_Array_10_21_reset = reset;
  assign PE_Array_10_21_io_in_activate = PE_Array_10_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_21_io_in_weight = PE_Array_9_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_21_io_in_psum = PE_Array_9_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_22_clock = clock;
  assign PE_Array_10_22_reset = reset;
  assign PE_Array_10_22_io_in_activate = PE_Array_10_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_22_io_in_weight = PE_Array_9_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_22_io_in_psum = PE_Array_9_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_23_clock = clock;
  assign PE_Array_10_23_reset = reset;
  assign PE_Array_10_23_io_in_activate = PE_Array_10_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_23_io_in_weight = PE_Array_9_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_23_io_in_psum = PE_Array_9_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_24_clock = clock;
  assign PE_Array_10_24_reset = reset;
  assign PE_Array_10_24_io_in_activate = PE_Array_10_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_24_io_in_weight = PE_Array_9_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_24_io_in_psum = PE_Array_9_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_25_clock = clock;
  assign PE_Array_10_25_reset = reset;
  assign PE_Array_10_25_io_in_activate = PE_Array_10_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_25_io_in_weight = PE_Array_9_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_25_io_in_psum = PE_Array_9_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_26_clock = clock;
  assign PE_Array_10_26_reset = reset;
  assign PE_Array_10_26_io_in_activate = PE_Array_10_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_26_io_in_weight = PE_Array_9_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_26_io_in_psum = PE_Array_9_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_27_clock = clock;
  assign PE_Array_10_27_reset = reset;
  assign PE_Array_10_27_io_in_activate = PE_Array_10_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_27_io_in_weight = PE_Array_9_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_27_io_in_psum = PE_Array_9_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_28_clock = clock;
  assign PE_Array_10_28_reset = reset;
  assign PE_Array_10_28_io_in_activate = PE_Array_10_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_28_io_in_weight = PE_Array_9_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_28_io_in_psum = PE_Array_9_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_29_clock = clock;
  assign PE_Array_10_29_reset = reset;
  assign PE_Array_10_29_io_in_activate = PE_Array_10_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_29_io_in_weight = PE_Array_9_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_29_io_in_psum = PE_Array_9_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_30_clock = clock;
  assign PE_Array_10_30_reset = reset;
  assign PE_Array_10_30_io_in_activate = PE_Array_10_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_30_io_in_weight = PE_Array_9_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_30_io_in_psum = PE_Array_9_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_10_31_clock = clock;
  assign PE_Array_10_31_reset = reset;
  assign PE_Array_10_31_io_in_activate = PE_Array_10_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_10_31_io_in_weight = PE_Array_9_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_10_31_io_in_psum = PE_Array_9_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_10_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_10_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_0_clock = clock;
  assign PE_Array_11_0_reset = reset;
  assign PE_Array_11_0_io_in_activate = io_activate_11; // @[DataPath.scala 11:26]
  assign PE_Array_11_0_io_in_weight = PE_Array_10_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_0_io_in_psum = PE_Array_10_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_1_clock = clock;
  assign PE_Array_11_1_reset = reset;
  assign PE_Array_11_1_io_in_activate = PE_Array_11_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_1_io_in_weight = PE_Array_10_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_1_io_in_psum = PE_Array_10_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_2_clock = clock;
  assign PE_Array_11_2_reset = reset;
  assign PE_Array_11_2_io_in_activate = PE_Array_11_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_2_io_in_weight = PE_Array_10_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_2_io_in_psum = PE_Array_10_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_3_clock = clock;
  assign PE_Array_11_3_reset = reset;
  assign PE_Array_11_3_io_in_activate = PE_Array_11_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_3_io_in_weight = PE_Array_10_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_3_io_in_psum = PE_Array_10_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_4_clock = clock;
  assign PE_Array_11_4_reset = reset;
  assign PE_Array_11_4_io_in_activate = PE_Array_11_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_4_io_in_weight = PE_Array_10_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_4_io_in_psum = PE_Array_10_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_5_clock = clock;
  assign PE_Array_11_5_reset = reset;
  assign PE_Array_11_5_io_in_activate = PE_Array_11_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_5_io_in_weight = PE_Array_10_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_5_io_in_psum = PE_Array_10_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_6_clock = clock;
  assign PE_Array_11_6_reset = reset;
  assign PE_Array_11_6_io_in_activate = PE_Array_11_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_6_io_in_weight = PE_Array_10_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_6_io_in_psum = PE_Array_10_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_7_clock = clock;
  assign PE_Array_11_7_reset = reset;
  assign PE_Array_11_7_io_in_activate = PE_Array_11_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_7_io_in_weight = PE_Array_10_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_7_io_in_psum = PE_Array_10_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_8_clock = clock;
  assign PE_Array_11_8_reset = reset;
  assign PE_Array_11_8_io_in_activate = PE_Array_11_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_8_io_in_weight = PE_Array_10_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_8_io_in_psum = PE_Array_10_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_9_clock = clock;
  assign PE_Array_11_9_reset = reset;
  assign PE_Array_11_9_io_in_activate = PE_Array_11_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_9_io_in_weight = PE_Array_10_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_9_io_in_psum = PE_Array_10_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_10_clock = clock;
  assign PE_Array_11_10_reset = reset;
  assign PE_Array_11_10_io_in_activate = PE_Array_11_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_10_io_in_weight = PE_Array_10_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_10_io_in_psum = PE_Array_10_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_11_clock = clock;
  assign PE_Array_11_11_reset = reset;
  assign PE_Array_11_11_io_in_activate = PE_Array_11_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_11_io_in_weight = PE_Array_10_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_11_io_in_psum = PE_Array_10_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_12_clock = clock;
  assign PE_Array_11_12_reset = reset;
  assign PE_Array_11_12_io_in_activate = PE_Array_11_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_12_io_in_weight = PE_Array_10_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_12_io_in_psum = PE_Array_10_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_13_clock = clock;
  assign PE_Array_11_13_reset = reset;
  assign PE_Array_11_13_io_in_activate = PE_Array_11_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_13_io_in_weight = PE_Array_10_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_13_io_in_psum = PE_Array_10_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_14_clock = clock;
  assign PE_Array_11_14_reset = reset;
  assign PE_Array_11_14_io_in_activate = PE_Array_11_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_14_io_in_weight = PE_Array_10_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_14_io_in_psum = PE_Array_10_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_15_clock = clock;
  assign PE_Array_11_15_reset = reset;
  assign PE_Array_11_15_io_in_activate = PE_Array_11_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_15_io_in_weight = PE_Array_10_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_15_io_in_psum = PE_Array_10_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_16_clock = clock;
  assign PE_Array_11_16_reset = reset;
  assign PE_Array_11_16_io_in_activate = PE_Array_11_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_16_io_in_weight = PE_Array_10_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_16_io_in_psum = PE_Array_10_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_17_clock = clock;
  assign PE_Array_11_17_reset = reset;
  assign PE_Array_11_17_io_in_activate = PE_Array_11_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_17_io_in_weight = PE_Array_10_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_17_io_in_psum = PE_Array_10_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_18_clock = clock;
  assign PE_Array_11_18_reset = reset;
  assign PE_Array_11_18_io_in_activate = PE_Array_11_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_18_io_in_weight = PE_Array_10_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_18_io_in_psum = PE_Array_10_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_19_clock = clock;
  assign PE_Array_11_19_reset = reset;
  assign PE_Array_11_19_io_in_activate = PE_Array_11_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_19_io_in_weight = PE_Array_10_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_19_io_in_psum = PE_Array_10_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_20_clock = clock;
  assign PE_Array_11_20_reset = reset;
  assign PE_Array_11_20_io_in_activate = PE_Array_11_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_20_io_in_weight = PE_Array_10_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_20_io_in_psum = PE_Array_10_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_21_clock = clock;
  assign PE_Array_11_21_reset = reset;
  assign PE_Array_11_21_io_in_activate = PE_Array_11_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_21_io_in_weight = PE_Array_10_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_21_io_in_psum = PE_Array_10_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_22_clock = clock;
  assign PE_Array_11_22_reset = reset;
  assign PE_Array_11_22_io_in_activate = PE_Array_11_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_22_io_in_weight = PE_Array_10_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_22_io_in_psum = PE_Array_10_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_23_clock = clock;
  assign PE_Array_11_23_reset = reset;
  assign PE_Array_11_23_io_in_activate = PE_Array_11_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_23_io_in_weight = PE_Array_10_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_23_io_in_psum = PE_Array_10_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_24_clock = clock;
  assign PE_Array_11_24_reset = reset;
  assign PE_Array_11_24_io_in_activate = PE_Array_11_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_24_io_in_weight = PE_Array_10_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_24_io_in_psum = PE_Array_10_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_25_clock = clock;
  assign PE_Array_11_25_reset = reset;
  assign PE_Array_11_25_io_in_activate = PE_Array_11_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_25_io_in_weight = PE_Array_10_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_25_io_in_psum = PE_Array_10_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_26_clock = clock;
  assign PE_Array_11_26_reset = reset;
  assign PE_Array_11_26_io_in_activate = PE_Array_11_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_26_io_in_weight = PE_Array_10_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_26_io_in_psum = PE_Array_10_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_27_clock = clock;
  assign PE_Array_11_27_reset = reset;
  assign PE_Array_11_27_io_in_activate = PE_Array_11_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_27_io_in_weight = PE_Array_10_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_27_io_in_psum = PE_Array_10_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_28_clock = clock;
  assign PE_Array_11_28_reset = reset;
  assign PE_Array_11_28_io_in_activate = PE_Array_11_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_28_io_in_weight = PE_Array_10_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_28_io_in_psum = PE_Array_10_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_29_clock = clock;
  assign PE_Array_11_29_reset = reset;
  assign PE_Array_11_29_io_in_activate = PE_Array_11_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_29_io_in_weight = PE_Array_10_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_29_io_in_psum = PE_Array_10_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_30_clock = clock;
  assign PE_Array_11_30_reset = reset;
  assign PE_Array_11_30_io_in_activate = PE_Array_11_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_30_io_in_weight = PE_Array_10_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_30_io_in_psum = PE_Array_10_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_11_31_clock = clock;
  assign PE_Array_11_31_reset = reset;
  assign PE_Array_11_31_io_in_activate = PE_Array_11_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_11_31_io_in_weight = PE_Array_10_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_11_31_io_in_psum = PE_Array_10_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_11_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_11_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_0_clock = clock;
  assign PE_Array_12_0_reset = reset;
  assign PE_Array_12_0_io_in_activate = io_activate_12; // @[DataPath.scala 11:26]
  assign PE_Array_12_0_io_in_weight = PE_Array_11_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_0_io_in_psum = PE_Array_11_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_1_clock = clock;
  assign PE_Array_12_1_reset = reset;
  assign PE_Array_12_1_io_in_activate = PE_Array_12_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_1_io_in_weight = PE_Array_11_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_1_io_in_psum = PE_Array_11_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_2_clock = clock;
  assign PE_Array_12_2_reset = reset;
  assign PE_Array_12_2_io_in_activate = PE_Array_12_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_2_io_in_weight = PE_Array_11_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_2_io_in_psum = PE_Array_11_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_3_clock = clock;
  assign PE_Array_12_3_reset = reset;
  assign PE_Array_12_3_io_in_activate = PE_Array_12_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_3_io_in_weight = PE_Array_11_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_3_io_in_psum = PE_Array_11_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_4_clock = clock;
  assign PE_Array_12_4_reset = reset;
  assign PE_Array_12_4_io_in_activate = PE_Array_12_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_4_io_in_weight = PE_Array_11_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_4_io_in_psum = PE_Array_11_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_5_clock = clock;
  assign PE_Array_12_5_reset = reset;
  assign PE_Array_12_5_io_in_activate = PE_Array_12_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_5_io_in_weight = PE_Array_11_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_5_io_in_psum = PE_Array_11_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_6_clock = clock;
  assign PE_Array_12_6_reset = reset;
  assign PE_Array_12_6_io_in_activate = PE_Array_12_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_6_io_in_weight = PE_Array_11_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_6_io_in_psum = PE_Array_11_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_7_clock = clock;
  assign PE_Array_12_7_reset = reset;
  assign PE_Array_12_7_io_in_activate = PE_Array_12_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_7_io_in_weight = PE_Array_11_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_7_io_in_psum = PE_Array_11_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_8_clock = clock;
  assign PE_Array_12_8_reset = reset;
  assign PE_Array_12_8_io_in_activate = PE_Array_12_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_8_io_in_weight = PE_Array_11_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_8_io_in_psum = PE_Array_11_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_9_clock = clock;
  assign PE_Array_12_9_reset = reset;
  assign PE_Array_12_9_io_in_activate = PE_Array_12_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_9_io_in_weight = PE_Array_11_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_9_io_in_psum = PE_Array_11_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_10_clock = clock;
  assign PE_Array_12_10_reset = reset;
  assign PE_Array_12_10_io_in_activate = PE_Array_12_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_10_io_in_weight = PE_Array_11_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_10_io_in_psum = PE_Array_11_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_11_clock = clock;
  assign PE_Array_12_11_reset = reset;
  assign PE_Array_12_11_io_in_activate = PE_Array_12_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_11_io_in_weight = PE_Array_11_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_11_io_in_psum = PE_Array_11_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_12_clock = clock;
  assign PE_Array_12_12_reset = reset;
  assign PE_Array_12_12_io_in_activate = PE_Array_12_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_12_io_in_weight = PE_Array_11_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_12_io_in_psum = PE_Array_11_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_13_clock = clock;
  assign PE_Array_12_13_reset = reset;
  assign PE_Array_12_13_io_in_activate = PE_Array_12_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_13_io_in_weight = PE_Array_11_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_13_io_in_psum = PE_Array_11_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_14_clock = clock;
  assign PE_Array_12_14_reset = reset;
  assign PE_Array_12_14_io_in_activate = PE_Array_12_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_14_io_in_weight = PE_Array_11_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_14_io_in_psum = PE_Array_11_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_15_clock = clock;
  assign PE_Array_12_15_reset = reset;
  assign PE_Array_12_15_io_in_activate = PE_Array_12_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_15_io_in_weight = PE_Array_11_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_15_io_in_psum = PE_Array_11_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_16_clock = clock;
  assign PE_Array_12_16_reset = reset;
  assign PE_Array_12_16_io_in_activate = PE_Array_12_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_16_io_in_weight = PE_Array_11_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_16_io_in_psum = PE_Array_11_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_17_clock = clock;
  assign PE_Array_12_17_reset = reset;
  assign PE_Array_12_17_io_in_activate = PE_Array_12_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_17_io_in_weight = PE_Array_11_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_17_io_in_psum = PE_Array_11_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_18_clock = clock;
  assign PE_Array_12_18_reset = reset;
  assign PE_Array_12_18_io_in_activate = PE_Array_12_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_18_io_in_weight = PE_Array_11_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_18_io_in_psum = PE_Array_11_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_19_clock = clock;
  assign PE_Array_12_19_reset = reset;
  assign PE_Array_12_19_io_in_activate = PE_Array_12_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_19_io_in_weight = PE_Array_11_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_19_io_in_psum = PE_Array_11_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_20_clock = clock;
  assign PE_Array_12_20_reset = reset;
  assign PE_Array_12_20_io_in_activate = PE_Array_12_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_20_io_in_weight = PE_Array_11_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_20_io_in_psum = PE_Array_11_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_21_clock = clock;
  assign PE_Array_12_21_reset = reset;
  assign PE_Array_12_21_io_in_activate = PE_Array_12_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_21_io_in_weight = PE_Array_11_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_21_io_in_psum = PE_Array_11_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_22_clock = clock;
  assign PE_Array_12_22_reset = reset;
  assign PE_Array_12_22_io_in_activate = PE_Array_12_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_22_io_in_weight = PE_Array_11_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_22_io_in_psum = PE_Array_11_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_23_clock = clock;
  assign PE_Array_12_23_reset = reset;
  assign PE_Array_12_23_io_in_activate = PE_Array_12_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_23_io_in_weight = PE_Array_11_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_23_io_in_psum = PE_Array_11_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_24_clock = clock;
  assign PE_Array_12_24_reset = reset;
  assign PE_Array_12_24_io_in_activate = PE_Array_12_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_24_io_in_weight = PE_Array_11_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_24_io_in_psum = PE_Array_11_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_25_clock = clock;
  assign PE_Array_12_25_reset = reset;
  assign PE_Array_12_25_io_in_activate = PE_Array_12_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_25_io_in_weight = PE_Array_11_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_25_io_in_psum = PE_Array_11_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_26_clock = clock;
  assign PE_Array_12_26_reset = reset;
  assign PE_Array_12_26_io_in_activate = PE_Array_12_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_26_io_in_weight = PE_Array_11_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_26_io_in_psum = PE_Array_11_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_27_clock = clock;
  assign PE_Array_12_27_reset = reset;
  assign PE_Array_12_27_io_in_activate = PE_Array_12_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_27_io_in_weight = PE_Array_11_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_27_io_in_psum = PE_Array_11_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_28_clock = clock;
  assign PE_Array_12_28_reset = reset;
  assign PE_Array_12_28_io_in_activate = PE_Array_12_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_28_io_in_weight = PE_Array_11_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_28_io_in_psum = PE_Array_11_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_29_clock = clock;
  assign PE_Array_12_29_reset = reset;
  assign PE_Array_12_29_io_in_activate = PE_Array_12_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_29_io_in_weight = PE_Array_11_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_29_io_in_psum = PE_Array_11_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_30_clock = clock;
  assign PE_Array_12_30_reset = reset;
  assign PE_Array_12_30_io_in_activate = PE_Array_12_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_30_io_in_weight = PE_Array_11_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_30_io_in_psum = PE_Array_11_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_12_31_clock = clock;
  assign PE_Array_12_31_reset = reset;
  assign PE_Array_12_31_io_in_activate = PE_Array_12_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_12_31_io_in_weight = PE_Array_11_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_12_31_io_in_psum = PE_Array_11_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_12_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_12_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_0_clock = clock;
  assign PE_Array_13_0_reset = reset;
  assign PE_Array_13_0_io_in_activate = io_activate_13; // @[DataPath.scala 11:26]
  assign PE_Array_13_0_io_in_weight = PE_Array_12_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_0_io_in_psum = PE_Array_12_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_1_clock = clock;
  assign PE_Array_13_1_reset = reset;
  assign PE_Array_13_1_io_in_activate = PE_Array_13_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_1_io_in_weight = PE_Array_12_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_1_io_in_psum = PE_Array_12_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_2_clock = clock;
  assign PE_Array_13_2_reset = reset;
  assign PE_Array_13_2_io_in_activate = PE_Array_13_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_2_io_in_weight = PE_Array_12_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_2_io_in_psum = PE_Array_12_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_3_clock = clock;
  assign PE_Array_13_3_reset = reset;
  assign PE_Array_13_3_io_in_activate = PE_Array_13_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_3_io_in_weight = PE_Array_12_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_3_io_in_psum = PE_Array_12_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_4_clock = clock;
  assign PE_Array_13_4_reset = reset;
  assign PE_Array_13_4_io_in_activate = PE_Array_13_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_4_io_in_weight = PE_Array_12_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_4_io_in_psum = PE_Array_12_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_5_clock = clock;
  assign PE_Array_13_5_reset = reset;
  assign PE_Array_13_5_io_in_activate = PE_Array_13_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_5_io_in_weight = PE_Array_12_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_5_io_in_psum = PE_Array_12_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_6_clock = clock;
  assign PE_Array_13_6_reset = reset;
  assign PE_Array_13_6_io_in_activate = PE_Array_13_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_6_io_in_weight = PE_Array_12_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_6_io_in_psum = PE_Array_12_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_7_clock = clock;
  assign PE_Array_13_7_reset = reset;
  assign PE_Array_13_7_io_in_activate = PE_Array_13_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_7_io_in_weight = PE_Array_12_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_7_io_in_psum = PE_Array_12_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_8_clock = clock;
  assign PE_Array_13_8_reset = reset;
  assign PE_Array_13_8_io_in_activate = PE_Array_13_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_8_io_in_weight = PE_Array_12_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_8_io_in_psum = PE_Array_12_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_9_clock = clock;
  assign PE_Array_13_9_reset = reset;
  assign PE_Array_13_9_io_in_activate = PE_Array_13_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_9_io_in_weight = PE_Array_12_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_9_io_in_psum = PE_Array_12_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_10_clock = clock;
  assign PE_Array_13_10_reset = reset;
  assign PE_Array_13_10_io_in_activate = PE_Array_13_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_10_io_in_weight = PE_Array_12_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_10_io_in_psum = PE_Array_12_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_11_clock = clock;
  assign PE_Array_13_11_reset = reset;
  assign PE_Array_13_11_io_in_activate = PE_Array_13_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_11_io_in_weight = PE_Array_12_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_11_io_in_psum = PE_Array_12_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_12_clock = clock;
  assign PE_Array_13_12_reset = reset;
  assign PE_Array_13_12_io_in_activate = PE_Array_13_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_12_io_in_weight = PE_Array_12_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_12_io_in_psum = PE_Array_12_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_13_clock = clock;
  assign PE_Array_13_13_reset = reset;
  assign PE_Array_13_13_io_in_activate = PE_Array_13_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_13_io_in_weight = PE_Array_12_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_13_io_in_psum = PE_Array_12_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_14_clock = clock;
  assign PE_Array_13_14_reset = reset;
  assign PE_Array_13_14_io_in_activate = PE_Array_13_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_14_io_in_weight = PE_Array_12_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_14_io_in_psum = PE_Array_12_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_15_clock = clock;
  assign PE_Array_13_15_reset = reset;
  assign PE_Array_13_15_io_in_activate = PE_Array_13_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_15_io_in_weight = PE_Array_12_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_15_io_in_psum = PE_Array_12_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_16_clock = clock;
  assign PE_Array_13_16_reset = reset;
  assign PE_Array_13_16_io_in_activate = PE_Array_13_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_16_io_in_weight = PE_Array_12_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_16_io_in_psum = PE_Array_12_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_17_clock = clock;
  assign PE_Array_13_17_reset = reset;
  assign PE_Array_13_17_io_in_activate = PE_Array_13_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_17_io_in_weight = PE_Array_12_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_17_io_in_psum = PE_Array_12_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_18_clock = clock;
  assign PE_Array_13_18_reset = reset;
  assign PE_Array_13_18_io_in_activate = PE_Array_13_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_18_io_in_weight = PE_Array_12_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_18_io_in_psum = PE_Array_12_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_19_clock = clock;
  assign PE_Array_13_19_reset = reset;
  assign PE_Array_13_19_io_in_activate = PE_Array_13_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_19_io_in_weight = PE_Array_12_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_19_io_in_psum = PE_Array_12_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_20_clock = clock;
  assign PE_Array_13_20_reset = reset;
  assign PE_Array_13_20_io_in_activate = PE_Array_13_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_20_io_in_weight = PE_Array_12_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_20_io_in_psum = PE_Array_12_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_21_clock = clock;
  assign PE_Array_13_21_reset = reset;
  assign PE_Array_13_21_io_in_activate = PE_Array_13_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_21_io_in_weight = PE_Array_12_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_21_io_in_psum = PE_Array_12_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_22_clock = clock;
  assign PE_Array_13_22_reset = reset;
  assign PE_Array_13_22_io_in_activate = PE_Array_13_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_22_io_in_weight = PE_Array_12_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_22_io_in_psum = PE_Array_12_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_23_clock = clock;
  assign PE_Array_13_23_reset = reset;
  assign PE_Array_13_23_io_in_activate = PE_Array_13_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_23_io_in_weight = PE_Array_12_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_23_io_in_psum = PE_Array_12_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_24_clock = clock;
  assign PE_Array_13_24_reset = reset;
  assign PE_Array_13_24_io_in_activate = PE_Array_13_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_24_io_in_weight = PE_Array_12_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_24_io_in_psum = PE_Array_12_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_25_clock = clock;
  assign PE_Array_13_25_reset = reset;
  assign PE_Array_13_25_io_in_activate = PE_Array_13_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_25_io_in_weight = PE_Array_12_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_25_io_in_psum = PE_Array_12_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_26_clock = clock;
  assign PE_Array_13_26_reset = reset;
  assign PE_Array_13_26_io_in_activate = PE_Array_13_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_26_io_in_weight = PE_Array_12_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_26_io_in_psum = PE_Array_12_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_27_clock = clock;
  assign PE_Array_13_27_reset = reset;
  assign PE_Array_13_27_io_in_activate = PE_Array_13_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_27_io_in_weight = PE_Array_12_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_27_io_in_psum = PE_Array_12_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_28_clock = clock;
  assign PE_Array_13_28_reset = reset;
  assign PE_Array_13_28_io_in_activate = PE_Array_13_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_28_io_in_weight = PE_Array_12_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_28_io_in_psum = PE_Array_12_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_29_clock = clock;
  assign PE_Array_13_29_reset = reset;
  assign PE_Array_13_29_io_in_activate = PE_Array_13_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_29_io_in_weight = PE_Array_12_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_29_io_in_psum = PE_Array_12_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_30_clock = clock;
  assign PE_Array_13_30_reset = reset;
  assign PE_Array_13_30_io_in_activate = PE_Array_13_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_30_io_in_weight = PE_Array_12_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_30_io_in_psum = PE_Array_12_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_13_31_clock = clock;
  assign PE_Array_13_31_reset = reset;
  assign PE_Array_13_31_io_in_activate = PE_Array_13_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_13_31_io_in_weight = PE_Array_12_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_13_31_io_in_psum = PE_Array_12_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_13_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_13_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_0_clock = clock;
  assign PE_Array_14_0_reset = reset;
  assign PE_Array_14_0_io_in_activate = io_activate_14; // @[DataPath.scala 11:26]
  assign PE_Array_14_0_io_in_weight = PE_Array_13_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_0_io_in_psum = PE_Array_13_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_1_clock = clock;
  assign PE_Array_14_1_reset = reset;
  assign PE_Array_14_1_io_in_activate = PE_Array_14_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_1_io_in_weight = PE_Array_13_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_1_io_in_psum = PE_Array_13_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_2_clock = clock;
  assign PE_Array_14_2_reset = reset;
  assign PE_Array_14_2_io_in_activate = PE_Array_14_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_2_io_in_weight = PE_Array_13_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_2_io_in_psum = PE_Array_13_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_3_clock = clock;
  assign PE_Array_14_3_reset = reset;
  assign PE_Array_14_3_io_in_activate = PE_Array_14_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_3_io_in_weight = PE_Array_13_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_3_io_in_psum = PE_Array_13_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_4_clock = clock;
  assign PE_Array_14_4_reset = reset;
  assign PE_Array_14_4_io_in_activate = PE_Array_14_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_4_io_in_weight = PE_Array_13_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_4_io_in_psum = PE_Array_13_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_5_clock = clock;
  assign PE_Array_14_5_reset = reset;
  assign PE_Array_14_5_io_in_activate = PE_Array_14_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_5_io_in_weight = PE_Array_13_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_5_io_in_psum = PE_Array_13_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_6_clock = clock;
  assign PE_Array_14_6_reset = reset;
  assign PE_Array_14_6_io_in_activate = PE_Array_14_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_6_io_in_weight = PE_Array_13_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_6_io_in_psum = PE_Array_13_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_7_clock = clock;
  assign PE_Array_14_7_reset = reset;
  assign PE_Array_14_7_io_in_activate = PE_Array_14_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_7_io_in_weight = PE_Array_13_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_7_io_in_psum = PE_Array_13_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_8_clock = clock;
  assign PE_Array_14_8_reset = reset;
  assign PE_Array_14_8_io_in_activate = PE_Array_14_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_8_io_in_weight = PE_Array_13_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_8_io_in_psum = PE_Array_13_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_9_clock = clock;
  assign PE_Array_14_9_reset = reset;
  assign PE_Array_14_9_io_in_activate = PE_Array_14_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_9_io_in_weight = PE_Array_13_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_9_io_in_psum = PE_Array_13_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_10_clock = clock;
  assign PE_Array_14_10_reset = reset;
  assign PE_Array_14_10_io_in_activate = PE_Array_14_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_10_io_in_weight = PE_Array_13_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_10_io_in_psum = PE_Array_13_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_11_clock = clock;
  assign PE_Array_14_11_reset = reset;
  assign PE_Array_14_11_io_in_activate = PE_Array_14_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_11_io_in_weight = PE_Array_13_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_11_io_in_psum = PE_Array_13_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_12_clock = clock;
  assign PE_Array_14_12_reset = reset;
  assign PE_Array_14_12_io_in_activate = PE_Array_14_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_12_io_in_weight = PE_Array_13_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_12_io_in_psum = PE_Array_13_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_13_clock = clock;
  assign PE_Array_14_13_reset = reset;
  assign PE_Array_14_13_io_in_activate = PE_Array_14_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_13_io_in_weight = PE_Array_13_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_13_io_in_psum = PE_Array_13_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_14_clock = clock;
  assign PE_Array_14_14_reset = reset;
  assign PE_Array_14_14_io_in_activate = PE_Array_14_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_14_io_in_weight = PE_Array_13_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_14_io_in_psum = PE_Array_13_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_15_clock = clock;
  assign PE_Array_14_15_reset = reset;
  assign PE_Array_14_15_io_in_activate = PE_Array_14_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_15_io_in_weight = PE_Array_13_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_15_io_in_psum = PE_Array_13_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_16_clock = clock;
  assign PE_Array_14_16_reset = reset;
  assign PE_Array_14_16_io_in_activate = PE_Array_14_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_16_io_in_weight = PE_Array_13_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_16_io_in_psum = PE_Array_13_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_17_clock = clock;
  assign PE_Array_14_17_reset = reset;
  assign PE_Array_14_17_io_in_activate = PE_Array_14_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_17_io_in_weight = PE_Array_13_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_17_io_in_psum = PE_Array_13_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_18_clock = clock;
  assign PE_Array_14_18_reset = reset;
  assign PE_Array_14_18_io_in_activate = PE_Array_14_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_18_io_in_weight = PE_Array_13_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_18_io_in_psum = PE_Array_13_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_19_clock = clock;
  assign PE_Array_14_19_reset = reset;
  assign PE_Array_14_19_io_in_activate = PE_Array_14_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_19_io_in_weight = PE_Array_13_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_19_io_in_psum = PE_Array_13_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_20_clock = clock;
  assign PE_Array_14_20_reset = reset;
  assign PE_Array_14_20_io_in_activate = PE_Array_14_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_20_io_in_weight = PE_Array_13_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_20_io_in_psum = PE_Array_13_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_21_clock = clock;
  assign PE_Array_14_21_reset = reset;
  assign PE_Array_14_21_io_in_activate = PE_Array_14_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_21_io_in_weight = PE_Array_13_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_21_io_in_psum = PE_Array_13_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_22_clock = clock;
  assign PE_Array_14_22_reset = reset;
  assign PE_Array_14_22_io_in_activate = PE_Array_14_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_22_io_in_weight = PE_Array_13_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_22_io_in_psum = PE_Array_13_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_23_clock = clock;
  assign PE_Array_14_23_reset = reset;
  assign PE_Array_14_23_io_in_activate = PE_Array_14_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_23_io_in_weight = PE_Array_13_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_23_io_in_psum = PE_Array_13_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_24_clock = clock;
  assign PE_Array_14_24_reset = reset;
  assign PE_Array_14_24_io_in_activate = PE_Array_14_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_24_io_in_weight = PE_Array_13_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_24_io_in_psum = PE_Array_13_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_25_clock = clock;
  assign PE_Array_14_25_reset = reset;
  assign PE_Array_14_25_io_in_activate = PE_Array_14_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_25_io_in_weight = PE_Array_13_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_25_io_in_psum = PE_Array_13_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_26_clock = clock;
  assign PE_Array_14_26_reset = reset;
  assign PE_Array_14_26_io_in_activate = PE_Array_14_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_26_io_in_weight = PE_Array_13_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_26_io_in_psum = PE_Array_13_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_27_clock = clock;
  assign PE_Array_14_27_reset = reset;
  assign PE_Array_14_27_io_in_activate = PE_Array_14_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_27_io_in_weight = PE_Array_13_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_27_io_in_psum = PE_Array_13_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_28_clock = clock;
  assign PE_Array_14_28_reset = reset;
  assign PE_Array_14_28_io_in_activate = PE_Array_14_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_28_io_in_weight = PE_Array_13_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_28_io_in_psum = PE_Array_13_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_29_clock = clock;
  assign PE_Array_14_29_reset = reset;
  assign PE_Array_14_29_io_in_activate = PE_Array_14_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_29_io_in_weight = PE_Array_13_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_29_io_in_psum = PE_Array_13_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_30_clock = clock;
  assign PE_Array_14_30_reset = reset;
  assign PE_Array_14_30_io_in_activate = PE_Array_14_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_30_io_in_weight = PE_Array_13_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_30_io_in_psum = PE_Array_13_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_14_31_clock = clock;
  assign PE_Array_14_31_reset = reset;
  assign PE_Array_14_31_io_in_activate = PE_Array_14_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_14_31_io_in_weight = PE_Array_13_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_14_31_io_in_psum = PE_Array_13_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_14_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_14_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_0_clock = clock;
  assign PE_Array_15_0_reset = reset;
  assign PE_Array_15_0_io_in_activate = io_activate_15; // @[DataPath.scala 11:26]
  assign PE_Array_15_0_io_in_weight = PE_Array_14_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_0_io_in_psum = PE_Array_14_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_1_clock = clock;
  assign PE_Array_15_1_reset = reset;
  assign PE_Array_15_1_io_in_activate = PE_Array_15_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_1_io_in_weight = PE_Array_14_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_1_io_in_psum = PE_Array_14_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_2_clock = clock;
  assign PE_Array_15_2_reset = reset;
  assign PE_Array_15_2_io_in_activate = PE_Array_15_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_2_io_in_weight = PE_Array_14_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_2_io_in_psum = PE_Array_14_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_3_clock = clock;
  assign PE_Array_15_3_reset = reset;
  assign PE_Array_15_3_io_in_activate = PE_Array_15_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_3_io_in_weight = PE_Array_14_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_3_io_in_psum = PE_Array_14_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_4_clock = clock;
  assign PE_Array_15_4_reset = reset;
  assign PE_Array_15_4_io_in_activate = PE_Array_15_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_4_io_in_weight = PE_Array_14_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_4_io_in_psum = PE_Array_14_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_5_clock = clock;
  assign PE_Array_15_5_reset = reset;
  assign PE_Array_15_5_io_in_activate = PE_Array_15_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_5_io_in_weight = PE_Array_14_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_5_io_in_psum = PE_Array_14_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_6_clock = clock;
  assign PE_Array_15_6_reset = reset;
  assign PE_Array_15_6_io_in_activate = PE_Array_15_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_6_io_in_weight = PE_Array_14_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_6_io_in_psum = PE_Array_14_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_7_clock = clock;
  assign PE_Array_15_7_reset = reset;
  assign PE_Array_15_7_io_in_activate = PE_Array_15_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_7_io_in_weight = PE_Array_14_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_7_io_in_psum = PE_Array_14_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_8_clock = clock;
  assign PE_Array_15_8_reset = reset;
  assign PE_Array_15_8_io_in_activate = PE_Array_15_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_8_io_in_weight = PE_Array_14_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_8_io_in_psum = PE_Array_14_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_9_clock = clock;
  assign PE_Array_15_9_reset = reset;
  assign PE_Array_15_9_io_in_activate = PE_Array_15_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_9_io_in_weight = PE_Array_14_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_9_io_in_psum = PE_Array_14_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_10_clock = clock;
  assign PE_Array_15_10_reset = reset;
  assign PE_Array_15_10_io_in_activate = PE_Array_15_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_10_io_in_weight = PE_Array_14_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_10_io_in_psum = PE_Array_14_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_11_clock = clock;
  assign PE_Array_15_11_reset = reset;
  assign PE_Array_15_11_io_in_activate = PE_Array_15_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_11_io_in_weight = PE_Array_14_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_11_io_in_psum = PE_Array_14_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_12_clock = clock;
  assign PE_Array_15_12_reset = reset;
  assign PE_Array_15_12_io_in_activate = PE_Array_15_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_12_io_in_weight = PE_Array_14_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_12_io_in_psum = PE_Array_14_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_13_clock = clock;
  assign PE_Array_15_13_reset = reset;
  assign PE_Array_15_13_io_in_activate = PE_Array_15_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_13_io_in_weight = PE_Array_14_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_13_io_in_psum = PE_Array_14_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_14_clock = clock;
  assign PE_Array_15_14_reset = reset;
  assign PE_Array_15_14_io_in_activate = PE_Array_15_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_14_io_in_weight = PE_Array_14_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_14_io_in_psum = PE_Array_14_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_15_clock = clock;
  assign PE_Array_15_15_reset = reset;
  assign PE_Array_15_15_io_in_activate = PE_Array_15_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_15_io_in_weight = PE_Array_14_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_15_io_in_psum = PE_Array_14_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_16_clock = clock;
  assign PE_Array_15_16_reset = reset;
  assign PE_Array_15_16_io_in_activate = PE_Array_15_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_16_io_in_weight = PE_Array_14_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_16_io_in_psum = PE_Array_14_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_17_clock = clock;
  assign PE_Array_15_17_reset = reset;
  assign PE_Array_15_17_io_in_activate = PE_Array_15_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_17_io_in_weight = PE_Array_14_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_17_io_in_psum = PE_Array_14_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_18_clock = clock;
  assign PE_Array_15_18_reset = reset;
  assign PE_Array_15_18_io_in_activate = PE_Array_15_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_18_io_in_weight = PE_Array_14_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_18_io_in_psum = PE_Array_14_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_19_clock = clock;
  assign PE_Array_15_19_reset = reset;
  assign PE_Array_15_19_io_in_activate = PE_Array_15_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_19_io_in_weight = PE_Array_14_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_19_io_in_psum = PE_Array_14_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_20_clock = clock;
  assign PE_Array_15_20_reset = reset;
  assign PE_Array_15_20_io_in_activate = PE_Array_15_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_20_io_in_weight = PE_Array_14_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_20_io_in_psum = PE_Array_14_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_21_clock = clock;
  assign PE_Array_15_21_reset = reset;
  assign PE_Array_15_21_io_in_activate = PE_Array_15_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_21_io_in_weight = PE_Array_14_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_21_io_in_psum = PE_Array_14_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_22_clock = clock;
  assign PE_Array_15_22_reset = reset;
  assign PE_Array_15_22_io_in_activate = PE_Array_15_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_22_io_in_weight = PE_Array_14_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_22_io_in_psum = PE_Array_14_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_23_clock = clock;
  assign PE_Array_15_23_reset = reset;
  assign PE_Array_15_23_io_in_activate = PE_Array_15_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_23_io_in_weight = PE_Array_14_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_23_io_in_psum = PE_Array_14_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_24_clock = clock;
  assign PE_Array_15_24_reset = reset;
  assign PE_Array_15_24_io_in_activate = PE_Array_15_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_24_io_in_weight = PE_Array_14_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_24_io_in_psum = PE_Array_14_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_25_clock = clock;
  assign PE_Array_15_25_reset = reset;
  assign PE_Array_15_25_io_in_activate = PE_Array_15_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_25_io_in_weight = PE_Array_14_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_25_io_in_psum = PE_Array_14_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_26_clock = clock;
  assign PE_Array_15_26_reset = reset;
  assign PE_Array_15_26_io_in_activate = PE_Array_15_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_26_io_in_weight = PE_Array_14_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_26_io_in_psum = PE_Array_14_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_27_clock = clock;
  assign PE_Array_15_27_reset = reset;
  assign PE_Array_15_27_io_in_activate = PE_Array_15_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_27_io_in_weight = PE_Array_14_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_27_io_in_psum = PE_Array_14_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_28_clock = clock;
  assign PE_Array_15_28_reset = reset;
  assign PE_Array_15_28_io_in_activate = PE_Array_15_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_28_io_in_weight = PE_Array_14_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_28_io_in_psum = PE_Array_14_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_29_clock = clock;
  assign PE_Array_15_29_reset = reset;
  assign PE_Array_15_29_io_in_activate = PE_Array_15_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_29_io_in_weight = PE_Array_14_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_29_io_in_psum = PE_Array_14_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_30_clock = clock;
  assign PE_Array_15_30_reset = reset;
  assign PE_Array_15_30_io_in_activate = PE_Array_15_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_30_io_in_weight = PE_Array_14_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_30_io_in_psum = PE_Array_14_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_15_31_clock = clock;
  assign PE_Array_15_31_reset = reset;
  assign PE_Array_15_31_io_in_activate = PE_Array_15_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_15_31_io_in_weight = PE_Array_14_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_15_31_io_in_psum = PE_Array_14_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_15_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_15_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_0_clock = clock;
  assign PE_Array_16_0_reset = reset;
  assign PE_Array_16_0_io_in_activate = io_activate_16; // @[DataPath.scala 11:26]
  assign PE_Array_16_0_io_in_weight = PE_Array_15_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_0_io_in_psum = PE_Array_15_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_1_clock = clock;
  assign PE_Array_16_1_reset = reset;
  assign PE_Array_16_1_io_in_activate = PE_Array_16_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_1_io_in_weight = PE_Array_15_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_1_io_in_psum = PE_Array_15_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_2_clock = clock;
  assign PE_Array_16_2_reset = reset;
  assign PE_Array_16_2_io_in_activate = PE_Array_16_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_2_io_in_weight = PE_Array_15_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_2_io_in_psum = PE_Array_15_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_3_clock = clock;
  assign PE_Array_16_3_reset = reset;
  assign PE_Array_16_3_io_in_activate = PE_Array_16_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_3_io_in_weight = PE_Array_15_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_3_io_in_psum = PE_Array_15_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_4_clock = clock;
  assign PE_Array_16_4_reset = reset;
  assign PE_Array_16_4_io_in_activate = PE_Array_16_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_4_io_in_weight = PE_Array_15_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_4_io_in_psum = PE_Array_15_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_5_clock = clock;
  assign PE_Array_16_5_reset = reset;
  assign PE_Array_16_5_io_in_activate = PE_Array_16_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_5_io_in_weight = PE_Array_15_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_5_io_in_psum = PE_Array_15_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_6_clock = clock;
  assign PE_Array_16_6_reset = reset;
  assign PE_Array_16_6_io_in_activate = PE_Array_16_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_6_io_in_weight = PE_Array_15_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_6_io_in_psum = PE_Array_15_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_7_clock = clock;
  assign PE_Array_16_7_reset = reset;
  assign PE_Array_16_7_io_in_activate = PE_Array_16_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_7_io_in_weight = PE_Array_15_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_7_io_in_psum = PE_Array_15_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_8_clock = clock;
  assign PE_Array_16_8_reset = reset;
  assign PE_Array_16_8_io_in_activate = PE_Array_16_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_8_io_in_weight = PE_Array_15_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_8_io_in_psum = PE_Array_15_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_9_clock = clock;
  assign PE_Array_16_9_reset = reset;
  assign PE_Array_16_9_io_in_activate = PE_Array_16_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_9_io_in_weight = PE_Array_15_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_9_io_in_psum = PE_Array_15_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_10_clock = clock;
  assign PE_Array_16_10_reset = reset;
  assign PE_Array_16_10_io_in_activate = PE_Array_16_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_10_io_in_weight = PE_Array_15_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_10_io_in_psum = PE_Array_15_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_11_clock = clock;
  assign PE_Array_16_11_reset = reset;
  assign PE_Array_16_11_io_in_activate = PE_Array_16_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_11_io_in_weight = PE_Array_15_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_11_io_in_psum = PE_Array_15_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_12_clock = clock;
  assign PE_Array_16_12_reset = reset;
  assign PE_Array_16_12_io_in_activate = PE_Array_16_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_12_io_in_weight = PE_Array_15_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_12_io_in_psum = PE_Array_15_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_13_clock = clock;
  assign PE_Array_16_13_reset = reset;
  assign PE_Array_16_13_io_in_activate = PE_Array_16_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_13_io_in_weight = PE_Array_15_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_13_io_in_psum = PE_Array_15_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_14_clock = clock;
  assign PE_Array_16_14_reset = reset;
  assign PE_Array_16_14_io_in_activate = PE_Array_16_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_14_io_in_weight = PE_Array_15_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_14_io_in_psum = PE_Array_15_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_15_clock = clock;
  assign PE_Array_16_15_reset = reset;
  assign PE_Array_16_15_io_in_activate = PE_Array_16_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_15_io_in_weight = PE_Array_15_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_15_io_in_psum = PE_Array_15_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_16_clock = clock;
  assign PE_Array_16_16_reset = reset;
  assign PE_Array_16_16_io_in_activate = PE_Array_16_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_16_io_in_weight = PE_Array_15_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_16_io_in_psum = PE_Array_15_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_17_clock = clock;
  assign PE_Array_16_17_reset = reset;
  assign PE_Array_16_17_io_in_activate = PE_Array_16_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_17_io_in_weight = PE_Array_15_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_17_io_in_psum = PE_Array_15_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_18_clock = clock;
  assign PE_Array_16_18_reset = reset;
  assign PE_Array_16_18_io_in_activate = PE_Array_16_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_18_io_in_weight = PE_Array_15_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_18_io_in_psum = PE_Array_15_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_19_clock = clock;
  assign PE_Array_16_19_reset = reset;
  assign PE_Array_16_19_io_in_activate = PE_Array_16_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_19_io_in_weight = PE_Array_15_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_19_io_in_psum = PE_Array_15_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_20_clock = clock;
  assign PE_Array_16_20_reset = reset;
  assign PE_Array_16_20_io_in_activate = PE_Array_16_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_20_io_in_weight = PE_Array_15_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_20_io_in_psum = PE_Array_15_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_21_clock = clock;
  assign PE_Array_16_21_reset = reset;
  assign PE_Array_16_21_io_in_activate = PE_Array_16_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_21_io_in_weight = PE_Array_15_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_21_io_in_psum = PE_Array_15_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_22_clock = clock;
  assign PE_Array_16_22_reset = reset;
  assign PE_Array_16_22_io_in_activate = PE_Array_16_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_22_io_in_weight = PE_Array_15_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_22_io_in_psum = PE_Array_15_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_23_clock = clock;
  assign PE_Array_16_23_reset = reset;
  assign PE_Array_16_23_io_in_activate = PE_Array_16_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_23_io_in_weight = PE_Array_15_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_23_io_in_psum = PE_Array_15_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_24_clock = clock;
  assign PE_Array_16_24_reset = reset;
  assign PE_Array_16_24_io_in_activate = PE_Array_16_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_24_io_in_weight = PE_Array_15_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_24_io_in_psum = PE_Array_15_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_25_clock = clock;
  assign PE_Array_16_25_reset = reset;
  assign PE_Array_16_25_io_in_activate = PE_Array_16_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_25_io_in_weight = PE_Array_15_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_25_io_in_psum = PE_Array_15_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_26_clock = clock;
  assign PE_Array_16_26_reset = reset;
  assign PE_Array_16_26_io_in_activate = PE_Array_16_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_26_io_in_weight = PE_Array_15_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_26_io_in_psum = PE_Array_15_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_27_clock = clock;
  assign PE_Array_16_27_reset = reset;
  assign PE_Array_16_27_io_in_activate = PE_Array_16_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_27_io_in_weight = PE_Array_15_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_27_io_in_psum = PE_Array_15_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_28_clock = clock;
  assign PE_Array_16_28_reset = reset;
  assign PE_Array_16_28_io_in_activate = PE_Array_16_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_28_io_in_weight = PE_Array_15_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_28_io_in_psum = PE_Array_15_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_29_clock = clock;
  assign PE_Array_16_29_reset = reset;
  assign PE_Array_16_29_io_in_activate = PE_Array_16_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_29_io_in_weight = PE_Array_15_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_29_io_in_psum = PE_Array_15_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_30_clock = clock;
  assign PE_Array_16_30_reset = reset;
  assign PE_Array_16_30_io_in_activate = PE_Array_16_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_30_io_in_weight = PE_Array_15_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_30_io_in_psum = PE_Array_15_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_16_31_clock = clock;
  assign PE_Array_16_31_reset = reset;
  assign PE_Array_16_31_io_in_activate = PE_Array_16_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_16_31_io_in_weight = PE_Array_15_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_16_31_io_in_psum = PE_Array_15_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_16_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_16_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_0_clock = clock;
  assign PE_Array_17_0_reset = reset;
  assign PE_Array_17_0_io_in_activate = io_activate_17; // @[DataPath.scala 11:26]
  assign PE_Array_17_0_io_in_weight = PE_Array_16_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_0_io_in_psum = PE_Array_16_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_1_clock = clock;
  assign PE_Array_17_1_reset = reset;
  assign PE_Array_17_1_io_in_activate = PE_Array_17_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_1_io_in_weight = PE_Array_16_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_1_io_in_psum = PE_Array_16_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_2_clock = clock;
  assign PE_Array_17_2_reset = reset;
  assign PE_Array_17_2_io_in_activate = PE_Array_17_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_2_io_in_weight = PE_Array_16_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_2_io_in_psum = PE_Array_16_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_3_clock = clock;
  assign PE_Array_17_3_reset = reset;
  assign PE_Array_17_3_io_in_activate = PE_Array_17_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_3_io_in_weight = PE_Array_16_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_3_io_in_psum = PE_Array_16_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_4_clock = clock;
  assign PE_Array_17_4_reset = reset;
  assign PE_Array_17_4_io_in_activate = PE_Array_17_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_4_io_in_weight = PE_Array_16_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_4_io_in_psum = PE_Array_16_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_5_clock = clock;
  assign PE_Array_17_5_reset = reset;
  assign PE_Array_17_5_io_in_activate = PE_Array_17_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_5_io_in_weight = PE_Array_16_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_5_io_in_psum = PE_Array_16_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_6_clock = clock;
  assign PE_Array_17_6_reset = reset;
  assign PE_Array_17_6_io_in_activate = PE_Array_17_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_6_io_in_weight = PE_Array_16_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_6_io_in_psum = PE_Array_16_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_7_clock = clock;
  assign PE_Array_17_7_reset = reset;
  assign PE_Array_17_7_io_in_activate = PE_Array_17_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_7_io_in_weight = PE_Array_16_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_7_io_in_psum = PE_Array_16_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_8_clock = clock;
  assign PE_Array_17_8_reset = reset;
  assign PE_Array_17_8_io_in_activate = PE_Array_17_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_8_io_in_weight = PE_Array_16_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_8_io_in_psum = PE_Array_16_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_9_clock = clock;
  assign PE_Array_17_9_reset = reset;
  assign PE_Array_17_9_io_in_activate = PE_Array_17_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_9_io_in_weight = PE_Array_16_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_9_io_in_psum = PE_Array_16_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_10_clock = clock;
  assign PE_Array_17_10_reset = reset;
  assign PE_Array_17_10_io_in_activate = PE_Array_17_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_10_io_in_weight = PE_Array_16_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_10_io_in_psum = PE_Array_16_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_11_clock = clock;
  assign PE_Array_17_11_reset = reset;
  assign PE_Array_17_11_io_in_activate = PE_Array_17_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_11_io_in_weight = PE_Array_16_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_11_io_in_psum = PE_Array_16_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_12_clock = clock;
  assign PE_Array_17_12_reset = reset;
  assign PE_Array_17_12_io_in_activate = PE_Array_17_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_12_io_in_weight = PE_Array_16_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_12_io_in_psum = PE_Array_16_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_13_clock = clock;
  assign PE_Array_17_13_reset = reset;
  assign PE_Array_17_13_io_in_activate = PE_Array_17_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_13_io_in_weight = PE_Array_16_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_13_io_in_psum = PE_Array_16_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_14_clock = clock;
  assign PE_Array_17_14_reset = reset;
  assign PE_Array_17_14_io_in_activate = PE_Array_17_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_14_io_in_weight = PE_Array_16_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_14_io_in_psum = PE_Array_16_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_15_clock = clock;
  assign PE_Array_17_15_reset = reset;
  assign PE_Array_17_15_io_in_activate = PE_Array_17_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_15_io_in_weight = PE_Array_16_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_15_io_in_psum = PE_Array_16_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_16_clock = clock;
  assign PE_Array_17_16_reset = reset;
  assign PE_Array_17_16_io_in_activate = PE_Array_17_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_16_io_in_weight = PE_Array_16_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_16_io_in_psum = PE_Array_16_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_17_clock = clock;
  assign PE_Array_17_17_reset = reset;
  assign PE_Array_17_17_io_in_activate = PE_Array_17_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_17_io_in_weight = PE_Array_16_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_17_io_in_psum = PE_Array_16_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_18_clock = clock;
  assign PE_Array_17_18_reset = reset;
  assign PE_Array_17_18_io_in_activate = PE_Array_17_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_18_io_in_weight = PE_Array_16_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_18_io_in_psum = PE_Array_16_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_19_clock = clock;
  assign PE_Array_17_19_reset = reset;
  assign PE_Array_17_19_io_in_activate = PE_Array_17_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_19_io_in_weight = PE_Array_16_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_19_io_in_psum = PE_Array_16_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_20_clock = clock;
  assign PE_Array_17_20_reset = reset;
  assign PE_Array_17_20_io_in_activate = PE_Array_17_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_20_io_in_weight = PE_Array_16_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_20_io_in_psum = PE_Array_16_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_21_clock = clock;
  assign PE_Array_17_21_reset = reset;
  assign PE_Array_17_21_io_in_activate = PE_Array_17_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_21_io_in_weight = PE_Array_16_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_21_io_in_psum = PE_Array_16_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_22_clock = clock;
  assign PE_Array_17_22_reset = reset;
  assign PE_Array_17_22_io_in_activate = PE_Array_17_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_22_io_in_weight = PE_Array_16_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_22_io_in_psum = PE_Array_16_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_23_clock = clock;
  assign PE_Array_17_23_reset = reset;
  assign PE_Array_17_23_io_in_activate = PE_Array_17_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_23_io_in_weight = PE_Array_16_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_23_io_in_psum = PE_Array_16_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_24_clock = clock;
  assign PE_Array_17_24_reset = reset;
  assign PE_Array_17_24_io_in_activate = PE_Array_17_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_24_io_in_weight = PE_Array_16_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_24_io_in_psum = PE_Array_16_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_25_clock = clock;
  assign PE_Array_17_25_reset = reset;
  assign PE_Array_17_25_io_in_activate = PE_Array_17_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_25_io_in_weight = PE_Array_16_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_25_io_in_psum = PE_Array_16_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_26_clock = clock;
  assign PE_Array_17_26_reset = reset;
  assign PE_Array_17_26_io_in_activate = PE_Array_17_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_26_io_in_weight = PE_Array_16_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_26_io_in_psum = PE_Array_16_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_27_clock = clock;
  assign PE_Array_17_27_reset = reset;
  assign PE_Array_17_27_io_in_activate = PE_Array_17_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_27_io_in_weight = PE_Array_16_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_27_io_in_psum = PE_Array_16_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_28_clock = clock;
  assign PE_Array_17_28_reset = reset;
  assign PE_Array_17_28_io_in_activate = PE_Array_17_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_28_io_in_weight = PE_Array_16_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_28_io_in_psum = PE_Array_16_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_29_clock = clock;
  assign PE_Array_17_29_reset = reset;
  assign PE_Array_17_29_io_in_activate = PE_Array_17_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_29_io_in_weight = PE_Array_16_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_29_io_in_psum = PE_Array_16_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_30_clock = clock;
  assign PE_Array_17_30_reset = reset;
  assign PE_Array_17_30_io_in_activate = PE_Array_17_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_30_io_in_weight = PE_Array_16_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_30_io_in_psum = PE_Array_16_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_17_31_clock = clock;
  assign PE_Array_17_31_reset = reset;
  assign PE_Array_17_31_io_in_activate = PE_Array_17_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_17_31_io_in_weight = PE_Array_16_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_17_31_io_in_psum = PE_Array_16_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_17_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_17_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_0_clock = clock;
  assign PE_Array_18_0_reset = reset;
  assign PE_Array_18_0_io_in_activate = io_activate_18; // @[DataPath.scala 11:26]
  assign PE_Array_18_0_io_in_weight = PE_Array_17_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_0_io_in_psum = PE_Array_17_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_1_clock = clock;
  assign PE_Array_18_1_reset = reset;
  assign PE_Array_18_1_io_in_activate = PE_Array_18_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_1_io_in_weight = PE_Array_17_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_1_io_in_psum = PE_Array_17_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_2_clock = clock;
  assign PE_Array_18_2_reset = reset;
  assign PE_Array_18_2_io_in_activate = PE_Array_18_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_2_io_in_weight = PE_Array_17_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_2_io_in_psum = PE_Array_17_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_3_clock = clock;
  assign PE_Array_18_3_reset = reset;
  assign PE_Array_18_3_io_in_activate = PE_Array_18_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_3_io_in_weight = PE_Array_17_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_3_io_in_psum = PE_Array_17_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_4_clock = clock;
  assign PE_Array_18_4_reset = reset;
  assign PE_Array_18_4_io_in_activate = PE_Array_18_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_4_io_in_weight = PE_Array_17_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_4_io_in_psum = PE_Array_17_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_5_clock = clock;
  assign PE_Array_18_5_reset = reset;
  assign PE_Array_18_5_io_in_activate = PE_Array_18_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_5_io_in_weight = PE_Array_17_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_5_io_in_psum = PE_Array_17_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_6_clock = clock;
  assign PE_Array_18_6_reset = reset;
  assign PE_Array_18_6_io_in_activate = PE_Array_18_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_6_io_in_weight = PE_Array_17_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_6_io_in_psum = PE_Array_17_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_7_clock = clock;
  assign PE_Array_18_7_reset = reset;
  assign PE_Array_18_7_io_in_activate = PE_Array_18_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_7_io_in_weight = PE_Array_17_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_7_io_in_psum = PE_Array_17_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_8_clock = clock;
  assign PE_Array_18_8_reset = reset;
  assign PE_Array_18_8_io_in_activate = PE_Array_18_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_8_io_in_weight = PE_Array_17_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_8_io_in_psum = PE_Array_17_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_9_clock = clock;
  assign PE_Array_18_9_reset = reset;
  assign PE_Array_18_9_io_in_activate = PE_Array_18_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_9_io_in_weight = PE_Array_17_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_9_io_in_psum = PE_Array_17_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_10_clock = clock;
  assign PE_Array_18_10_reset = reset;
  assign PE_Array_18_10_io_in_activate = PE_Array_18_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_10_io_in_weight = PE_Array_17_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_10_io_in_psum = PE_Array_17_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_11_clock = clock;
  assign PE_Array_18_11_reset = reset;
  assign PE_Array_18_11_io_in_activate = PE_Array_18_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_11_io_in_weight = PE_Array_17_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_11_io_in_psum = PE_Array_17_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_12_clock = clock;
  assign PE_Array_18_12_reset = reset;
  assign PE_Array_18_12_io_in_activate = PE_Array_18_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_12_io_in_weight = PE_Array_17_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_12_io_in_psum = PE_Array_17_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_13_clock = clock;
  assign PE_Array_18_13_reset = reset;
  assign PE_Array_18_13_io_in_activate = PE_Array_18_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_13_io_in_weight = PE_Array_17_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_13_io_in_psum = PE_Array_17_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_14_clock = clock;
  assign PE_Array_18_14_reset = reset;
  assign PE_Array_18_14_io_in_activate = PE_Array_18_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_14_io_in_weight = PE_Array_17_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_14_io_in_psum = PE_Array_17_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_15_clock = clock;
  assign PE_Array_18_15_reset = reset;
  assign PE_Array_18_15_io_in_activate = PE_Array_18_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_15_io_in_weight = PE_Array_17_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_15_io_in_psum = PE_Array_17_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_16_clock = clock;
  assign PE_Array_18_16_reset = reset;
  assign PE_Array_18_16_io_in_activate = PE_Array_18_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_16_io_in_weight = PE_Array_17_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_16_io_in_psum = PE_Array_17_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_17_clock = clock;
  assign PE_Array_18_17_reset = reset;
  assign PE_Array_18_17_io_in_activate = PE_Array_18_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_17_io_in_weight = PE_Array_17_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_17_io_in_psum = PE_Array_17_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_18_clock = clock;
  assign PE_Array_18_18_reset = reset;
  assign PE_Array_18_18_io_in_activate = PE_Array_18_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_18_io_in_weight = PE_Array_17_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_18_io_in_psum = PE_Array_17_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_19_clock = clock;
  assign PE_Array_18_19_reset = reset;
  assign PE_Array_18_19_io_in_activate = PE_Array_18_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_19_io_in_weight = PE_Array_17_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_19_io_in_psum = PE_Array_17_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_20_clock = clock;
  assign PE_Array_18_20_reset = reset;
  assign PE_Array_18_20_io_in_activate = PE_Array_18_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_20_io_in_weight = PE_Array_17_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_20_io_in_psum = PE_Array_17_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_21_clock = clock;
  assign PE_Array_18_21_reset = reset;
  assign PE_Array_18_21_io_in_activate = PE_Array_18_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_21_io_in_weight = PE_Array_17_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_21_io_in_psum = PE_Array_17_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_22_clock = clock;
  assign PE_Array_18_22_reset = reset;
  assign PE_Array_18_22_io_in_activate = PE_Array_18_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_22_io_in_weight = PE_Array_17_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_22_io_in_psum = PE_Array_17_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_23_clock = clock;
  assign PE_Array_18_23_reset = reset;
  assign PE_Array_18_23_io_in_activate = PE_Array_18_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_23_io_in_weight = PE_Array_17_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_23_io_in_psum = PE_Array_17_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_24_clock = clock;
  assign PE_Array_18_24_reset = reset;
  assign PE_Array_18_24_io_in_activate = PE_Array_18_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_24_io_in_weight = PE_Array_17_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_24_io_in_psum = PE_Array_17_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_25_clock = clock;
  assign PE_Array_18_25_reset = reset;
  assign PE_Array_18_25_io_in_activate = PE_Array_18_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_25_io_in_weight = PE_Array_17_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_25_io_in_psum = PE_Array_17_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_26_clock = clock;
  assign PE_Array_18_26_reset = reset;
  assign PE_Array_18_26_io_in_activate = PE_Array_18_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_26_io_in_weight = PE_Array_17_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_26_io_in_psum = PE_Array_17_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_27_clock = clock;
  assign PE_Array_18_27_reset = reset;
  assign PE_Array_18_27_io_in_activate = PE_Array_18_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_27_io_in_weight = PE_Array_17_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_27_io_in_psum = PE_Array_17_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_28_clock = clock;
  assign PE_Array_18_28_reset = reset;
  assign PE_Array_18_28_io_in_activate = PE_Array_18_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_28_io_in_weight = PE_Array_17_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_28_io_in_psum = PE_Array_17_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_29_clock = clock;
  assign PE_Array_18_29_reset = reset;
  assign PE_Array_18_29_io_in_activate = PE_Array_18_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_29_io_in_weight = PE_Array_17_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_29_io_in_psum = PE_Array_17_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_30_clock = clock;
  assign PE_Array_18_30_reset = reset;
  assign PE_Array_18_30_io_in_activate = PE_Array_18_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_30_io_in_weight = PE_Array_17_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_30_io_in_psum = PE_Array_17_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_18_31_clock = clock;
  assign PE_Array_18_31_reset = reset;
  assign PE_Array_18_31_io_in_activate = PE_Array_18_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_18_31_io_in_weight = PE_Array_17_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_18_31_io_in_psum = PE_Array_17_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_18_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_18_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_0_clock = clock;
  assign PE_Array_19_0_reset = reset;
  assign PE_Array_19_0_io_in_activate = io_activate_19; // @[DataPath.scala 11:26]
  assign PE_Array_19_0_io_in_weight = PE_Array_18_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_0_io_in_psum = PE_Array_18_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_1_clock = clock;
  assign PE_Array_19_1_reset = reset;
  assign PE_Array_19_1_io_in_activate = PE_Array_19_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_1_io_in_weight = PE_Array_18_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_1_io_in_psum = PE_Array_18_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_2_clock = clock;
  assign PE_Array_19_2_reset = reset;
  assign PE_Array_19_2_io_in_activate = PE_Array_19_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_2_io_in_weight = PE_Array_18_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_2_io_in_psum = PE_Array_18_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_3_clock = clock;
  assign PE_Array_19_3_reset = reset;
  assign PE_Array_19_3_io_in_activate = PE_Array_19_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_3_io_in_weight = PE_Array_18_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_3_io_in_psum = PE_Array_18_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_4_clock = clock;
  assign PE_Array_19_4_reset = reset;
  assign PE_Array_19_4_io_in_activate = PE_Array_19_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_4_io_in_weight = PE_Array_18_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_4_io_in_psum = PE_Array_18_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_5_clock = clock;
  assign PE_Array_19_5_reset = reset;
  assign PE_Array_19_5_io_in_activate = PE_Array_19_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_5_io_in_weight = PE_Array_18_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_5_io_in_psum = PE_Array_18_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_6_clock = clock;
  assign PE_Array_19_6_reset = reset;
  assign PE_Array_19_6_io_in_activate = PE_Array_19_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_6_io_in_weight = PE_Array_18_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_6_io_in_psum = PE_Array_18_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_7_clock = clock;
  assign PE_Array_19_7_reset = reset;
  assign PE_Array_19_7_io_in_activate = PE_Array_19_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_7_io_in_weight = PE_Array_18_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_7_io_in_psum = PE_Array_18_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_8_clock = clock;
  assign PE_Array_19_8_reset = reset;
  assign PE_Array_19_8_io_in_activate = PE_Array_19_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_8_io_in_weight = PE_Array_18_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_8_io_in_psum = PE_Array_18_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_9_clock = clock;
  assign PE_Array_19_9_reset = reset;
  assign PE_Array_19_9_io_in_activate = PE_Array_19_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_9_io_in_weight = PE_Array_18_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_9_io_in_psum = PE_Array_18_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_10_clock = clock;
  assign PE_Array_19_10_reset = reset;
  assign PE_Array_19_10_io_in_activate = PE_Array_19_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_10_io_in_weight = PE_Array_18_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_10_io_in_psum = PE_Array_18_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_11_clock = clock;
  assign PE_Array_19_11_reset = reset;
  assign PE_Array_19_11_io_in_activate = PE_Array_19_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_11_io_in_weight = PE_Array_18_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_11_io_in_psum = PE_Array_18_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_12_clock = clock;
  assign PE_Array_19_12_reset = reset;
  assign PE_Array_19_12_io_in_activate = PE_Array_19_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_12_io_in_weight = PE_Array_18_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_12_io_in_psum = PE_Array_18_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_13_clock = clock;
  assign PE_Array_19_13_reset = reset;
  assign PE_Array_19_13_io_in_activate = PE_Array_19_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_13_io_in_weight = PE_Array_18_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_13_io_in_psum = PE_Array_18_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_14_clock = clock;
  assign PE_Array_19_14_reset = reset;
  assign PE_Array_19_14_io_in_activate = PE_Array_19_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_14_io_in_weight = PE_Array_18_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_14_io_in_psum = PE_Array_18_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_15_clock = clock;
  assign PE_Array_19_15_reset = reset;
  assign PE_Array_19_15_io_in_activate = PE_Array_19_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_15_io_in_weight = PE_Array_18_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_15_io_in_psum = PE_Array_18_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_16_clock = clock;
  assign PE_Array_19_16_reset = reset;
  assign PE_Array_19_16_io_in_activate = PE_Array_19_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_16_io_in_weight = PE_Array_18_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_16_io_in_psum = PE_Array_18_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_17_clock = clock;
  assign PE_Array_19_17_reset = reset;
  assign PE_Array_19_17_io_in_activate = PE_Array_19_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_17_io_in_weight = PE_Array_18_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_17_io_in_psum = PE_Array_18_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_18_clock = clock;
  assign PE_Array_19_18_reset = reset;
  assign PE_Array_19_18_io_in_activate = PE_Array_19_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_18_io_in_weight = PE_Array_18_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_18_io_in_psum = PE_Array_18_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_19_clock = clock;
  assign PE_Array_19_19_reset = reset;
  assign PE_Array_19_19_io_in_activate = PE_Array_19_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_19_io_in_weight = PE_Array_18_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_19_io_in_psum = PE_Array_18_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_20_clock = clock;
  assign PE_Array_19_20_reset = reset;
  assign PE_Array_19_20_io_in_activate = PE_Array_19_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_20_io_in_weight = PE_Array_18_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_20_io_in_psum = PE_Array_18_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_21_clock = clock;
  assign PE_Array_19_21_reset = reset;
  assign PE_Array_19_21_io_in_activate = PE_Array_19_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_21_io_in_weight = PE_Array_18_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_21_io_in_psum = PE_Array_18_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_22_clock = clock;
  assign PE_Array_19_22_reset = reset;
  assign PE_Array_19_22_io_in_activate = PE_Array_19_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_22_io_in_weight = PE_Array_18_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_22_io_in_psum = PE_Array_18_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_23_clock = clock;
  assign PE_Array_19_23_reset = reset;
  assign PE_Array_19_23_io_in_activate = PE_Array_19_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_23_io_in_weight = PE_Array_18_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_23_io_in_psum = PE_Array_18_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_24_clock = clock;
  assign PE_Array_19_24_reset = reset;
  assign PE_Array_19_24_io_in_activate = PE_Array_19_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_24_io_in_weight = PE_Array_18_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_24_io_in_psum = PE_Array_18_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_25_clock = clock;
  assign PE_Array_19_25_reset = reset;
  assign PE_Array_19_25_io_in_activate = PE_Array_19_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_25_io_in_weight = PE_Array_18_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_25_io_in_psum = PE_Array_18_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_26_clock = clock;
  assign PE_Array_19_26_reset = reset;
  assign PE_Array_19_26_io_in_activate = PE_Array_19_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_26_io_in_weight = PE_Array_18_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_26_io_in_psum = PE_Array_18_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_27_clock = clock;
  assign PE_Array_19_27_reset = reset;
  assign PE_Array_19_27_io_in_activate = PE_Array_19_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_27_io_in_weight = PE_Array_18_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_27_io_in_psum = PE_Array_18_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_28_clock = clock;
  assign PE_Array_19_28_reset = reset;
  assign PE_Array_19_28_io_in_activate = PE_Array_19_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_28_io_in_weight = PE_Array_18_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_28_io_in_psum = PE_Array_18_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_29_clock = clock;
  assign PE_Array_19_29_reset = reset;
  assign PE_Array_19_29_io_in_activate = PE_Array_19_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_29_io_in_weight = PE_Array_18_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_29_io_in_psum = PE_Array_18_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_30_clock = clock;
  assign PE_Array_19_30_reset = reset;
  assign PE_Array_19_30_io_in_activate = PE_Array_19_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_30_io_in_weight = PE_Array_18_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_30_io_in_psum = PE_Array_18_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_19_31_clock = clock;
  assign PE_Array_19_31_reset = reset;
  assign PE_Array_19_31_io_in_activate = PE_Array_19_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_19_31_io_in_weight = PE_Array_18_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_19_31_io_in_psum = PE_Array_18_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_19_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_19_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_0_clock = clock;
  assign PE_Array_20_0_reset = reset;
  assign PE_Array_20_0_io_in_activate = io_activate_20; // @[DataPath.scala 11:26]
  assign PE_Array_20_0_io_in_weight = PE_Array_19_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_0_io_in_psum = PE_Array_19_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_1_clock = clock;
  assign PE_Array_20_1_reset = reset;
  assign PE_Array_20_1_io_in_activate = PE_Array_20_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_1_io_in_weight = PE_Array_19_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_1_io_in_psum = PE_Array_19_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_2_clock = clock;
  assign PE_Array_20_2_reset = reset;
  assign PE_Array_20_2_io_in_activate = PE_Array_20_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_2_io_in_weight = PE_Array_19_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_2_io_in_psum = PE_Array_19_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_3_clock = clock;
  assign PE_Array_20_3_reset = reset;
  assign PE_Array_20_3_io_in_activate = PE_Array_20_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_3_io_in_weight = PE_Array_19_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_3_io_in_psum = PE_Array_19_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_4_clock = clock;
  assign PE_Array_20_4_reset = reset;
  assign PE_Array_20_4_io_in_activate = PE_Array_20_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_4_io_in_weight = PE_Array_19_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_4_io_in_psum = PE_Array_19_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_5_clock = clock;
  assign PE_Array_20_5_reset = reset;
  assign PE_Array_20_5_io_in_activate = PE_Array_20_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_5_io_in_weight = PE_Array_19_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_5_io_in_psum = PE_Array_19_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_6_clock = clock;
  assign PE_Array_20_6_reset = reset;
  assign PE_Array_20_6_io_in_activate = PE_Array_20_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_6_io_in_weight = PE_Array_19_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_6_io_in_psum = PE_Array_19_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_7_clock = clock;
  assign PE_Array_20_7_reset = reset;
  assign PE_Array_20_7_io_in_activate = PE_Array_20_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_7_io_in_weight = PE_Array_19_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_7_io_in_psum = PE_Array_19_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_8_clock = clock;
  assign PE_Array_20_8_reset = reset;
  assign PE_Array_20_8_io_in_activate = PE_Array_20_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_8_io_in_weight = PE_Array_19_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_8_io_in_psum = PE_Array_19_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_9_clock = clock;
  assign PE_Array_20_9_reset = reset;
  assign PE_Array_20_9_io_in_activate = PE_Array_20_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_9_io_in_weight = PE_Array_19_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_9_io_in_psum = PE_Array_19_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_10_clock = clock;
  assign PE_Array_20_10_reset = reset;
  assign PE_Array_20_10_io_in_activate = PE_Array_20_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_10_io_in_weight = PE_Array_19_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_10_io_in_psum = PE_Array_19_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_11_clock = clock;
  assign PE_Array_20_11_reset = reset;
  assign PE_Array_20_11_io_in_activate = PE_Array_20_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_11_io_in_weight = PE_Array_19_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_11_io_in_psum = PE_Array_19_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_12_clock = clock;
  assign PE_Array_20_12_reset = reset;
  assign PE_Array_20_12_io_in_activate = PE_Array_20_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_12_io_in_weight = PE_Array_19_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_12_io_in_psum = PE_Array_19_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_13_clock = clock;
  assign PE_Array_20_13_reset = reset;
  assign PE_Array_20_13_io_in_activate = PE_Array_20_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_13_io_in_weight = PE_Array_19_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_13_io_in_psum = PE_Array_19_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_14_clock = clock;
  assign PE_Array_20_14_reset = reset;
  assign PE_Array_20_14_io_in_activate = PE_Array_20_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_14_io_in_weight = PE_Array_19_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_14_io_in_psum = PE_Array_19_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_15_clock = clock;
  assign PE_Array_20_15_reset = reset;
  assign PE_Array_20_15_io_in_activate = PE_Array_20_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_15_io_in_weight = PE_Array_19_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_15_io_in_psum = PE_Array_19_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_16_clock = clock;
  assign PE_Array_20_16_reset = reset;
  assign PE_Array_20_16_io_in_activate = PE_Array_20_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_16_io_in_weight = PE_Array_19_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_16_io_in_psum = PE_Array_19_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_17_clock = clock;
  assign PE_Array_20_17_reset = reset;
  assign PE_Array_20_17_io_in_activate = PE_Array_20_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_17_io_in_weight = PE_Array_19_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_17_io_in_psum = PE_Array_19_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_18_clock = clock;
  assign PE_Array_20_18_reset = reset;
  assign PE_Array_20_18_io_in_activate = PE_Array_20_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_18_io_in_weight = PE_Array_19_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_18_io_in_psum = PE_Array_19_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_19_clock = clock;
  assign PE_Array_20_19_reset = reset;
  assign PE_Array_20_19_io_in_activate = PE_Array_20_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_19_io_in_weight = PE_Array_19_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_19_io_in_psum = PE_Array_19_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_20_clock = clock;
  assign PE_Array_20_20_reset = reset;
  assign PE_Array_20_20_io_in_activate = PE_Array_20_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_20_io_in_weight = PE_Array_19_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_20_io_in_psum = PE_Array_19_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_21_clock = clock;
  assign PE_Array_20_21_reset = reset;
  assign PE_Array_20_21_io_in_activate = PE_Array_20_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_21_io_in_weight = PE_Array_19_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_21_io_in_psum = PE_Array_19_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_22_clock = clock;
  assign PE_Array_20_22_reset = reset;
  assign PE_Array_20_22_io_in_activate = PE_Array_20_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_22_io_in_weight = PE_Array_19_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_22_io_in_psum = PE_Array_19_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_23_clock = clock;
  assign PE_Array_20_23_reset = reset;
  assign PE_Array_20_23_io_in_activate = PE_Array_20_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_23_io_in_weight = PE_Array_19_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_23_io_in_psum = PE_Array_19_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_24_clock = clock;
  assign PE_Array_20_24_reset = reset;
  assign PE_Array_20_24_io_in_activate = PE_Array_20_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_24_io_in_weight = PE_Array_19_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_24_io_in_psum = PE_Array_19_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_25_clock = clock;
  assign PE_Array_20_25_reset = reset;
  assign PE_Array_20_25_io_in_activate = PE_Array_20_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_25_io_in_weight = PE_Array_19_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_25_io_in_psum = PE_Array_19_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_26_clock = clock;
  assign PE_Array_20_26_reset = reset;
  assign PE_Array_20_26_io_in_activate = PE_Array_20_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_26_io_in_weight = PE_Array_19_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_26_io_in_psum = PE_Array_19_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_27_clock = clock;
  assign PE_Array_20_27_reset = reset;
  assign PE_Array_20_27_io_in_activate = PE_Array_20_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_27_io_in_weight = PE_Array_19_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_27_io_in_psum = PE_Array_19_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_28_clock = clock;
  assign PE_Array_20_28_reset = reset;
  assign PE_Array_20_28_io_in_activate = PE_Array_20_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_28_io_in_weight = PE_Array_19_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_28_io_in_psum = PE_Array_19_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_29_clock = clock;
  assign PE_Array_20_29_reset = reset;
  assign PE_Array_20_29_io_in_activate = PE_Array_20_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_29_io_in_weight = PE_Array_19_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_29_io_in_psum = PE_Array_19_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_30_clock = clock;
  assign PE_Array_20_30_reset = reset;
  assign PE_Array_20_30_io_in_activate = PE_Array_20_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_30_io_in_weight = PE_Array_19_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_30_io_in_psum = PE_Array_19_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_20_31_clock = clock;
  assign PE_Array_20_31_reset = reset;
  assign PE_Array_20_31_io_in_activate = PE_Array_20_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_20_31_io_in_weight = PE_Array_19_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_20_31_io_in_psum = PE_Array_19_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_20_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_20_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_0_clock = clock;
  assign PE_Array_21_0_reset = reset;
  assign PE_Array_21_0_io_in_activate = io_activate_21; // @[DataPath.scala 11:26]
  assign PE_Array_21_0_io_in_weight = PE_Array_20_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_0_io_in_psum = PE_Array_20_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_1_clock = clock;
  assign PE_Array_21_1_reset = reset;
  assign PE_Array_21_1_io_in_activate = PE_Array_21_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_1_io_in_weight = PE_Array_20_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_1_io_in_psum = PE_Array_20_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_2_clock = clock;
  assign PE_Array_21_2_reset = reset;
  assign PE_Array_21_2_io_in_activate = PE_Array_21_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_2_io_in_weight = PE_Array_20_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_2_io_in_psum = PE_Array_20_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_3_clock = clock;
  assign PE_Array_21_3_reset = reset;
  assign PE_Array_21_3_io_in_activate = PE_Array_21_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_3_io_in_weight = PE_Array_20_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_3_io_in_psum = PE_Array_20_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_4_clock = clock;
  assign PE_Array_21_4_reset = reset;
  assign PE_Array_21_4_io_in_activate = PE_Array_21_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_4_io_in_weight = PE_Array_20_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_4_io_in_psum = PE_Array_20_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_5_clock = clock;
  assign PE_Array_21_5_reset = reset;
  assign PE_Array_21_5_io_in_activate = PE_Array_21_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_5_io_in_weight = PE_Array_20_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_5_io_in_psum = PE_Array_20_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_6_clock = clock;
  assign PE_Array_21_6_reset = reset;
  assign PE_Array_21_6_io_in_activate = PE_Array_21_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_6_io_in_weight = PE_Array_20_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_6_io_in_psum = PE_Array_20_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_7_clock = clock;
  assign PE_Array_21_7_reset = reset;
  assign PE_Array_21_7_io_in_activate = PE_Array_21_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_7_io_in_weight = PE_Array_20_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_7_io_in_psum = PE_Array_20_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_8_clock = clock;
  assign PE_Array_21_8_reset = reset;
  assign PE_Array_21_8_io_in_activate = PE_Array_21_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_8_io_in_weight = PE_Array_20_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_8_io_in_psum = PE_Array_20_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_9_clock = clock;
  assign PE_Array_21_9_reset = reset;
  assign PE_Array_21_9_io_in_activate = PE_Array_21_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_9_io_in_weight = PE_Array_20_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_9_io_in_psum = PE_Array_20_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_10_clock = clock;
  assign PE_Array_21_10_reset = reset;
  assign PE_Array_21_10_io_in_activate = PE_Array_21_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_10_io_in_weight = PE_Array_20_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_10_io_in_psum = PE_Array_20_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_11_clock = clock;
  assign PE_Array_21_11_reset = reset;
  assign PE_Array_21_11_io_in_activate = PE_Array_21_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_11_io_in_weight = PE_Array_20_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_11_io_in_psum = PE_Array_20_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_12_clock = clock;
  assign PE_Array_21_12_reset = reset;
  assign PE_Array_21_12_io_in_activate = PE_Array_21_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_12_io_in_weight = PE_Array_20_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_12_io_in_psum = PE_Array_20_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_13_clock = clock;
  assign PE_Array_21_13_reset = reset;
  assign PE_Array_21_13_io_in_activate = PE_Array_21_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_13_io_in_weight = PE_Array_20_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_13_io_in_psum = PE_Array_20_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_14_clock = clock;
  assign PE_Array_21_14_reset = reset;
  assign PE_Array_21_14_io_in_activate = PE_Array_21_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_14_io_in_weight = PE_Array_20_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_14_io_in_psum = PE_Array_20_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_15_clock = clock;
  assign PE_Array_21_15_reset = reset;
  assign PE_Array_21_15_io_in_activate = PE_Array_21_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_15_io_in_weight = PE_Array_20_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_15_io_in_psum = PE_Array_20_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_16_clock = clock;
  assign PE_Array_21_16_reset = reset;
  assign PE_Array_21_16_io_in_activate = PE_Array_21_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_16_io_in_weight = PE_Array_20_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_16_io_in_psum = PE_Array_20_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_17_clock = clock;
  assign PE_Array_21_17_reset = reset;
  assign PE_Array_21_17_io_in_activate = PE_Array_21_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_17_io_in_weight = PE_Array_20_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_17_io_in_psum = PE_Array_20_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_18_clock = clock;
  assign PE_Array_21_18_reset = reset;
  assign PE_Array_21_18_io_in_activate = PE_Array_21_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_18_io_in_weight = PE_Array_20_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_18_io_in_psum = PE_Array_20_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_19_clock = clock;
  assign PE_Array_21_19_reset = reset;
  assign PE_Array_21_19_io_in_activate = PE_Array_21_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_19_io_in_weight = PE_Array_20_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_19_io_in_psum = PE_Array_20_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_20_clock = clock;
  assign PE_Array_21_20_reset = reset;
  assign PE_Array_21_20_io_in_activate = PE_Array_21_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_20_io_in_weight = PE_Array_20_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_20_io_in_psum = PE_Array_20_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_21_clock = clock;
  assign PE_Array_21_21_reset = reset;
  assign PE_Array_21_21_io_in_activate = PE_Array_21_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_21_io_in_weight = PE_Array_20_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_21_io_in_psum = PE_Array_20_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_22_clock = clock;
  assign PE_Array_21_22_reset = reset;
  assign PE_Array_21_22_io_in_activate = PE_Array_21_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_22_io_in_weight = PE_Array_20_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_22_io_in_psum = PE_Array_20_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_23_clock = clock;
  assign PE_Array_21_23_reset = reset;
  assign PE_Array_21_23_io_in_activate = PE_Array_21_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_23_io_in_weight = PE_Array_20_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_23_io_in_psum = PE_Array_20_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_24_clock = clock;
  assign PE_Array_21_24_reset = reset;
  assign PE_Array_21_24_io_in_activate = PE_Array_21_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_24_io_in_weight = PE_Array_20_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_24_io_in_psum = PE_Array_20_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_25_clock = clock;
  assign PE_Array_21_25_reset = reset;
  assign PE_Array_21_25_io_in_activate = PE_Array_21_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_25_io_in_weight = PE_Array_20_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_25_io_in_psum = PE_Array_20_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_26_clock = clock;
  assign PE_Array_21_26_reset = reset;
  assign PE_Array_21_26_io_in_activate = PE_Array_21_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_26_io_in_weight = PE_Array_20_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_26_io_in_psum = PE_Array_20_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_27_clock = clock;
  assign PE_Array_21_27_reset = reset;
  assign PE_Array_21_27_io_in_activate = PE_Array_21_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_27_io_in_weight = PE_Array_20_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_27_io_in_psum = PE_Array_20_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_28_clock = clock;
  assign PE_Array_21_28_reset = reset;
  assign PE_Array_21_28_io_in_activate = PE_Array_21_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_28_io_in_weight = PE_Array_20_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_28_io_in_psum = PE_Array_20_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_29_clock = clock;
  assign PE_Array_21_29_reset = reset;
  assign PE_Array_21_29_io_in_activate = PE_Array_21_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_29_io_in_weight = PE_Array_20_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_29_io_in_psum = PE_Array_20_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_30_clock = clock;
  assign PE_Array_21_30_reset = reset;
  assign PE_Array_21_30_io_in_activate = PE_Array_21_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_30_io_in_weight = PE_Array_20_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_30_io_in_psum = PE_Array_20_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_21_31_clock = clock;
  assign PE_Array_21_31_reset = reset;
  assign PE_Array_21_31_io_in_activate = PE_Array_21_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_21_31_io_in_weight = PE_Array_20_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_21_31_io_in_psum = PE_Array_20_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_21_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_21_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_0_clock = clock;
  assign PE_Array_22_0_reset = reset;
  assign PE_Array_22_0_io_in_activate = io_activate_22; // @[DataPath.scala 11:26]
  assign PE_Array_22_0_io_in_weight = PE_Array_21_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_0_io_in_psum = PE_Array_21_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_1_clock = clock;
  assign PE_Array_22_1_reset = reset;
  assign PE_Array_22_1_io_in_activate = PE_Array_22_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_1_io_in_weight = PE_Array_21_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_1_io_in_psum = PE_Array_21_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_2_clock = clock;
  assign PE_Array_22_2_reset = reset;
  assign PE_Array_22_2_io_in_activate = PE_Array_22_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_2_io_in_weight = PE_Array_21_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_2_io_in_psum = PE_Array_21_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_3_clock = clock;
  assign PE_Array_22_3_reset = reset;
  assign PE_Array_22_3_io_in_activate = PE_Array_22_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_3_io_in_weight = PE_Array_21_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_3_io_in_psum = PE_Array_21_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_4_clock = clock;
  assign PE_Array_22_4_reset = reset;
  assign PE_Array_22_4_io_in_activate = PE_Array_22_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_4_io_in_weight = PE_Array_21_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_4_io_in_psum = PE_Array_21_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_5_clock = clock;
  assign PE_Array_22_5_reset = reset;
  assign PE_Array_22_5_io_in_activate = PE_Array_22_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_5_io_in_weight = PE_Array_21_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_5_io_in_psum = PE_Array_21_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_6_clock = clock;
  assign PE_Array_22_6_reset = reset;
  assign PE_Array_22_6_io_in_activate = PE_Array_22_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_6_io_in_weight = PE_Array_21_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_6_io_in_psum = PE_Array_21_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_7_clock = clock;
  assign PE_Array_22_7_reset = reset;
  assign PE_Array_22_7_io_in_activate = PE_Array_22_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_7_io_in_weight = PE_Array_21_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_7_io_in_psum = PE_Array_21_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_8_clock = clock;
  assign PE_Array_22_8_reset = reset;
  assign PE_Array_22_8_io_in_activate = PE_Array_22_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_8_io_in_weight = PE_Array_21_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_8_io_in_psum = PE_Array_21_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_9_clock = clock;
  assign PE_Array_22_9_reset = reset;
  assign PE_Array_22_9_io_in_activate = PE_Array_22_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_9_io_in_weight = PE_Array_21_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_9_io_in_psum = PE_Array_21_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_10_clock = clock;
  assign PE_Array_22_10_reset = reset;
  assign PE_Array_22_10_io_in_activate = PE_Array_22_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_10_io_in_weight = PE_Array_21_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_10_io_in_psum = PE_Array_21_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_11_clock = clock;
  assign PE_Array_22_11_reset = reset;
  assign PE_Array_22_11_io_in_activate = PE_Array_22_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_11_io_in_weight = PE_Array_21_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_11_io_in_psum = PE_Array_21_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_12_clock = clock;
  assign PE_Array_22_12_reset = reset;
  assign PE_Array_22_12_io_in_activate = PE_Array_22_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_12_io_in_weight = PE_Array_21_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_12_io_in_psum = PE_Array_21_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_13_clock = clock;
  assign PE_Array_22_13_reset = reset;
  assign PE_Array_22_13_io_in_activate = PE_Array_22_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_13_io_in_weight = PE_Array_21_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_13_io_in_psum = PE_Array_21_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_14_clock = clock;
  assign PE_Array_22_14_reset = reset;
  assign PE_Array_22_14_io_in_activate = PE_Array_22_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_14_io_in_weight = PE_Array_21_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_14_io_in_psum = PE_Array_21_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_15_clock = clock;
  assign PE_Array_22_15_reset = reset;
  assign PE_Array_22_15_io_in_activate = PE_Array_22_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_15_io_in_weight = PE_Array_21_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_15_io_in_psum = PE_Array_21_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_16_clock = clock;
  assign PE_Array_22_16_reset = reset;
  assign PE_Array_22_16_io_in_activate = PE_Array_22_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_16_io_in_weight = PE_Array_21_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_16_io_in_psum = PE_Array_21_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_17_clock = clock;
  assign PE_Array_22_17_reset = reset;
  assign PE_Array_22_17_io_in_activate = PE_Array_22_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_17_io_in_weight = PE_Array_21_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_17_io_in_psum = PE_Array_21_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_18_clock = clock;
  assign PE_Array_22_18_reset = reset;
  assign PE_Array_22_18_io_in_activate = PE_Array_22_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_18_io_in_weight = PE_Array_21_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_18_io_in_psum = PE_Array_21_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_19_clock = clock;
  assign PE_Array_22_19_reset = reset;
  assign PE_Array_22_19_io_in_activate = PE_Array_22_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_19_io_in_weight = PE_Array_21_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_19_io_in_psum = PE_Array_21_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_20_clock = clock;
  assign PE_Array_22_20_reset = reset;
  assign PE_Array_22_20_io_in_activate = PE_Array_22_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_20_io_in_weight = PE_Array_21_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_20_io_in_psum = PE_Array_21_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_21_clock = clock;
  assign PE_Array_22_21_reset = reset;
  assign PE_Array_22_21_io_in_activate = PE_Array_22_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_21_io_in_weight = PE_Array_21_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_21_io_in_psum = PE_Array_21_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_22_clock = clock;
  assign PE_Array_22_22_reset = reset;
  assign PE_Array_22_22_io_in_activate = PE_Array_22_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_22_io_in_weight = PE_Array_21_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_22_io_in_psum = PE_Array_21_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_23_clock = clock;
  assign PE_Array_22_23_reset = reset;
  assign PE_Array_22_23_io_in_activate = PE_Array_22_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_23_io_in_weight = PE_Array_21_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_23_io_in_psum = PE_Array_21_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_24_clock = clock;
  assign PE_Array_22_24_reset = reset;
  assign PE_Array_22_24_io_in_activate = PE_Array_22_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_24_io_in_weight = PE_Array_21_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_24_io_in_psum = PE_Array_21_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_25_clock = clock;
  assign PE_Array_22_25_reset = reset;
  assign PE_Array_22_25_io_in_activate = PE_Array_22_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_25_io_in_weight = PE_Array_21_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_25_io_in_psum = PE_Array_21_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_26_clock = clock;
  assign PE_Array_22_26_reset = reset;
  assign PE_Array_22_26_io_in_activate = PE_Array_22_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_26_io_in_weight = PE_Array_21_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_26_io_in_psum = PE_Array_21_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_27_clock = clock;
  assign PE_Array_22_27_reset = reset;
  assign PE_Array_22_27_io_in_activate = PE_Array_22_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_27_io_in_weight = PE_Array_21_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_27_io_in_psum = PE_Array_21_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_28_clock = clock;
  assign PE_Array_22_28_reset = reset;
  assign PE_Array_22_28_io_in_activate = PE_Array_22_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_28_io_in_weight = PE_Array_21_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_28_io_in_psum = PE_Array_21_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_29_clock = clock;
  assign PE_Array_22_29_reset = reset;
  assign PE_Array_22_29_io_in_activate = PE_Array_22_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_29_io_in_weight = PE_Array_21_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_29_io_in_psum = PE_Array_21_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_30_clock = clock;
  assign PE_Array_22_30_reset = reset;
  assign PE_Array_22_30_io_in_activate = PE_Array_22_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_30_io_in_weight = PE_Array_21_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_30_io_in_psum = PE_Array_21_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_22_31_clock = clock;
  assign PE_Array_22_31_reset = reset;
  assign PE_Array_22_31_io_in_activate = PE_Array_22_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_22_31_io_in_weight = PE_Array_21_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_22_31_io_in_psum = PE_Array_21_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_22_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_22_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_0_clock = clock;
  assign PE_Array_23_0_reset = reset;
  assign PE_Array_23_0_io_in_activate = io_activate_23; // @[DataPath.scala 11:26]
  assign PE_Array_23_0_io_in_weight = PE_Array_22_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_0_io_in_psum = PE_Array_22_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_1_clock = clock;
  assign PE_Array_23_1_reset = reset;
  assign PE_Array_23_1_io_in_activate = PE_Array_23_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_1_io_in_weight = PE_Array_22_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_1_io_in_psum = PE_Array_22_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_2_clock = clock;
  assign PE_Array_23_2_reset = reset;
  assign PE_Array_23_2_io_in_activate = PE_Array_23_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_2_io_in_weight = PE_Array_22_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_2_io_in_psum = PE_Array_22_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_3_clock = clock;
  assign PE_Array_23_3_reset = reset;
  assign PE_Array_23_3_io_in_activate = PE_Array_23_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_3_io_in_weight = PE_Array_22_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_3_io_in_psum = PE_Array_22_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_4_clock = clock;
  assign PE_Array_23_4_reset = reset;
  assign PE_Array_23_4_io_in_activate = PE_Array_23_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_4_io_in_weight = PE_Array_22_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_4_io_in_psum = PE_Array_22_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_5_clock = clock;
  assign PE_Array_23_5_reset = reset;
  assign PE_Array_23_5_io_in_activate = PE_Array_23_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_5_io_in_weight = PE_Array_22_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_5_io_in_psum = PE_Array_22_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_6_clock = clock;
  assign PE_Array_23_6_reset = reset;
  assign PE_Array_23_6_io_in_activate = PE_Array_23_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_6_io_in_weight = PE_Array_22_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_6_io_in_psum = PE_Array_22_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_7_clock = clock;
  assign PE_Array_23_7_reset = reset;
  assign PE_Array_23_7_io_in_activate = PE_Array_23_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_7_io_in_weight = PE_Array_22_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_7_io_in_psum = PE_Array_22_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_8_clock = clock;
  assign PE_Array_23_8_reset = reset;
  assign PE_Array_23_8_io_in_activate = PE_Array_23_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_8_io_in_weight = PE_Array_22_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_8_io_in_psum = PE_Array_22_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_9_clock = clock;
  assign PE_Array_23_9_reset = reset;
  assign PE_Array_23_9_io_in_activate = PE_Array_23_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_9_io_in_weight = PE_Array_22_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_9_io_in_psum = PE_Array_22_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_10_clock = clock;
  assign PE_Array_23_10_reset = reset;
  assign PE_Array_23_10_io_in_activate = PE_Array_23_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_10_io_in_weight = PE_Array_22_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_10_io_in_psum = PE_Array_22_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_11_clock = clock;
  assign PE_Array_23_11_reset = reset;
  assign PE_Array_23_11_io_in_activate = PE_Array_23_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_11_io_in_weight = PE_Array_22_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_11_io_in_psum = PE_Array_22_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_12_clock = clock;
  assign PE_Array_23_12_reset = reset;
  assign PE_Array_23_12_io_in_activate = PE_Array_23_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_12_io_in_weight = PE_Array_22_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_12_io_in_psum = PE_Array_22_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_13_clock = clock;
  assign PE_Array_23_13_reset = reset;
  assign PE_Array_23_13_io_in_activate = PE_Array_23_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_13_io_in_weight = PE_Array_22_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_13_io_in_psum = PE_Array_22_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_14_clock = clock;
  assign PE_Array_23_14_reset = reset;
  assign PE_Array_23_14_io_in_activate = PE_Array_23_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_14_io_in_weight = PE_Array_22_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_14_io_in_psum = PE_Array_22_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_15_clock = clock;
  assign PE_Array_23_15_reset = reset;
  assign PE_Array_23_15_io_in_activate = PE_Array_23_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_15_io_in_weight = PE_Array_22_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_15_io_in_psum = PE_Array_22_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_16_clock = clock;
  assign PE_Array_23_16_reset = reset;
  assign PE_Array_23_16_io_in_activate = PE_Array_23_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_16_io_in_weight = PE_Array_22_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_16_io_in_psum = PE_Array_22_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_17_clock = clock;
  assign PE_Array_23_17_reset = reset;
  assign PE_Array_23_17_io_in_activate = PE_Array_23_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_17_io_in_weight = PE_Array_22_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_17_io_in_psum = PE_Array_22_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_18_clock = clock;
  assign PE_Array_23_18_reset = reset;
  assign PE_Array_23_18_io_in_activate = PE_Array_23_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_18_io_in_weight = PE_Array_22_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_18_io_in_psum = PE_Array_22_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_19_clock = clock;
  assign PE_Array_23_19_reset = reset;
  assign PE_Array_23_19_io_in_activate = PE_Array_23_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_19_io_in_weight = PE_Array_22_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_19_io_in_psum = PE_Array_22_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_20_clock = clock;
  assign PE_Array_23_20_reset = reset;
  assign PE_Array_23_20_io_in_activate = PE_Array_23_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_20_io_in_weight = PE_Array_22_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_20_io_in_psum = PE_Array_22_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_21_clock = clock;
  assign PE_Array_23_21_reset = reset;
  assign PE_Array_23_21_io_in_activate = PE_Array_23_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_21_io_in_weight = PE_Array_22_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_21_io_in_psum = PE_Array_22_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_22_clock = clock;
  assign PE_Array_23_22_reset = reset;
  assign PE_Array_23_22_io_in_activate = PE_Array_23_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_22_io_in_weight = PE_Array_22_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_22_io_in_psum = PE_Array_22_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_23_clock = clock;
  assign PE_Array_23_23_reset = reset;
  assign PE_Array_23_23_io_in_activate = PE_Array_23_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_23_io_in_weight = PE_Array_22_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_23_io_in_psum = PE_Array_22_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_24_clock = clock;
  assign PE_Array_23_24_reset = reset;
  assign PE_Array_23_24_io_in_activate = PE_Array_23_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_24_io_in_weight = PE_Array_22_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_24_io_in_psum = PE_Array_22_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_25_clock = clock;
  assign PE_Array_23_25_reset = reset;
  assign PE_Array_23_25_io_in_activate = PE_Array_23_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_25_io_in_weight = PE_Array_22_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_25_io_in_psum = PE_Array_22_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_26_clock = clock;
  assign PE_Array_23_26_reset = reset;
  assign PE_Array_23_26_io_in_activate = PE_Array_23_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_26_io_in_weight = PE_Array_22_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_26_io_in_psum = PE_Array_22_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_27_clock = clock;
  assign PE_Array_23_27_reset = reset;
  assign PE_Array_23_27_io_in_activate = PE_Array_23_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_27_io_in_weight = PE_Array_22_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_27_io_in_psum = PE_Array_22_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_28_clock = clock;
  assign PE_Array_23_28_reset = reset;
  assign PE_Array_23_28_io_in_activate = PE_Array_23_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_28_io_in_weight = PE_Array_22_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_28_io_in_psum = PE_Array_22_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_29_clock = clock;
  assign PE_Array_23_29_reset = reset;
  assign PE_Array_23_29_io_in_activate = PE_Array_23_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_29_io_in_weight = PE_Array_22_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_29_io_in_psum = PE_Array_22_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_30_clock = clock;
  assign PE_Array_23_30_reset = reset;
  assign PE_Array_23_30_io_in_activate = PE_Array_23_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_30_io_in_weight = PE_Array_22_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_30_io_in_psum = PE_Array_22_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_23_31_clock = clock;
  assign PE_Array_23_31_reset = reset;
  assign PE_Array_23_31_io_in_activate = PE_Array_23_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_23_31_io_in_weight = PE_Array_22_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_23_31_io_in_psum = PE_Array_22_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_23_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_23_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_0_clock = clock;
  assign PE_Array_24_0_reset = reset;
  assign PE_Array_24_0_io_in_activate = io_activate_24; // @[DataPath.scala 11:26]
  assign PE_Array_24_0_io_in_weight = PE_Array_23_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_0_io_in_psum = PE_Array_23_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_1_clock = clock;
  assign PE_Array_24_1_reset = reset;
  assign PE_Array_24_1_io_in_activate = PE_Array_24_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_1_io_in_weight = PE_Array_23_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_1_io_in_psum = PE_Array_23_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_2_clock = clock;
  assign PE_Array_24_2_reset = reset;
  assign PE_Array_24_2_io_in_activate = PE_Array_24_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_2_io_in_weight = PE_Array_23_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_2_io_in_psum = PE_Array_23_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_3_clock = clock;
  assign PE_Array_24_3_reset = reset;
  assign PE_Array_24_3_io_in_activate = PE_Array_24_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_3_io_in_weight = PE_Array_23_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_3_io_in_psum = PE_Array_23_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_4_clock = clock;
  assign PE_Array_24_4_reset = reset;
  assign PE_Array_24_4_io_in_activate = PE_Array_24_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_4_io_in_weight = PE_Array_23_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_4_io_in_psum = PE_Array_23_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_5_clock = clock;
  assign PE_Array_24_5_reset = reset;
  assign PE_Array_24_5_io_in_activate = PE_Array_24_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_5_io_in_weight = PE_Array_23_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_5_io_in_psum = PE_Array_23_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_6_clock = clock;
  assign PE_Array_24_6_reset = reset;
  assign PE_Array_24_6_io_in_activate = PE_Array_24_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_6_io_in_weight = PE_Array_23_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_6_io_in_psum = PE_Array_23_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_7_clock = clock;
  assign PE_Array_24_7_reset = reset;
  assign PE_Array_24_7_io_in_activate = PE_Array_24_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_7_io_in_weight = PE_Array_23_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_7_io_in_psum = PE_Array_23_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_8_clock = clock;
  assign PE_Array_24_8_reset = reset;
  assign PE_Array_24_8_io_in_activate = PE_Array_24_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_8_io_in_weight = PE_Array_23_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_8_io_in_psum = PE_Array_23_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_9_clock = clock;
  assign PE_Array_24_9_reset = reset;
  assign PE_Array_24_9_io_in_activate = PE_Array_24_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_9_io_in_weight = PE_Array_23_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_9_io_in_psum = PE_Array_23_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_10_clock = clock;
  assign PE_Array_24_10_reset = reset;
  assign PE_Array_24_10_io_in_activate = PE_Array_24_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_10_io_in_weight = PE_Array_23_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_10_io_in_psum = PE_Array_23_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_11_clock = clock;
  assign PE_Array_24_11_reset = reset;
  assign PE_Array_24_11_io_in_activate = PE_Array_24_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_11_io_in_weight = PE_Array_23_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_11_io_in_psum = PE_Array_23_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_12_clock = clock;
  assign PE_Array_24_12_reset = reset;
  assign PE_Array_24_12_io_in_activate = PE_Array_24_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_12_io_in_weight = PE_Array_23_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_12_io_in_psum = PE_Array_23_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_13_clock = clock;
  assign PE_Array_24_13_reset = reset;
  assign PE_Array_24_13_io_in_activate = PE_Array_24_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_13_io_in_weight = PE_Array_23_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_13_io_in_psum = PE_Array_23_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_14_clock = clock;
  assign PE_Array_24_14_reset = reset;
  assign PE_Array_24_14_io_in_activate = PE_Array_24_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_14_io_in_weight = PE_Array_23_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_14_io_in_psum = PE_Array_23_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_15_clock = clock;
  assign PE_Array_24_15_reset = reset;
  assign PE_Array_24_15_io_in_activate = PE_Array_24_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_15_io_in_weight = PE_Array_23_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_15_io_in_psum = PE_Array_23_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_16_clock = clock;
  assign PE_Array_24_16_reset = reset;
  assign PE_Array_24_16_io_in_activate = PE_Array_24_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_16_io_in_weight = PE_Array_23_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_16_io_in_psum = PE_Array_23_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_17_clock = clock;
  assign PE_Array_24_17_reset = reset;
  assign PE_Array_24_17_io_in_activate = PE_Array_24_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_17_io_in_weight = PE_Array_23_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_17_io_in_psum = PE_Array_23_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_18_clock = clock;
  assign PE_Array_24_18_reset = reset;
  assign PE_Array_24_18_io_in_activate = PE_Array_24_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_18_io_in_weight = PE_Array_23_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_18_io_in_psum = PE_Array_23_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_19_clock = clock;
  assign PE_Array_24_19_reset = reset;
  assign PE_Array_24_19_io_in_activate = PE_Array_24_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_19_io_in_weight = PE_Array_23_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_19_io_in_psum = PE_Array_23_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_20_clock = clock;
  assign PE_Array_24_20_reset = reset;
  assign PE_Array_24_20_io_in_activate = PE_Array_24_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_20_io_in_weight = PE_Array_23_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_20_io_in_psum = PE_Array_23_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_21_clock = clock;
  assign PE_Array_24_21_reset = reset;
  assign PE_Array_24_21_io_in_activate = PE_Array_24_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_21_io_in_weight = PE_Array_23_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_21_io_in_psum = PE_Array_23_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_22_clock = clock;
  assign PE_Array_24_22_reset = reset;
  assign PE_Array_24_22_io_in_activate = PE_Array_24_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_22_io_in_weight = PE_Array_23_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_22_io_in_psum = PE_Array_23_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_23_clock = clock;
  assign PE_Array_24_23_reset = reset;
  assign PE_Array_24_23_io_in_activate = PE_Array_24_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_23_io_in_weight = PE_Array_23_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_23_io_in_psum = PE_Array_23_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_24_clock = clock;
  assign PE_Array_24_24_reset = reset;
  assign PE_Array_24_24_io_in_activate = PE_Array_24_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_24_io_in_weight = PE_Array_23_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_24_io_in_psum = PE_Array_23_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_25_clock = clock;
  assign PE_Array_24_25_reset = reset;
  assign PE_Array_24_25_io_in_activate = PE_Array_24_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_25_io_in_weight = PE_Array_23_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_25_io_in_psum = PE_Array_23_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_26_clock = clock;
  assign PE_Array_24_26_reset = reset;
  assign PE_Array_24_26_io_in_activate = PE_Array_24_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_26_io_in_weight = PE_Array_23_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_26_io_in_psum = PE_Array_23_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_27_clock = clock;
  assign PE_Array_24_27_reset = reset;
  assign PE_Array_24_27_io_in_activate = PE_Array_24_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_27_io_in_weight = PE_Array_23_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_27_io_in_psum = PE_Array_23_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_28_clock = clock;
  assign PE_Array_24_28_reset = reset;
  assign PE_Array_24_28_io_in_activate = PE_Array_24_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_28_io_in_weight = PE_Array_23_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_28_io_in_psum = PE_Array_23_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_29_clock = clock;
  assign PE_Array_24_29_reset = reset;
  assign PE_Array_24_29_io_in_activate = PE_Array_24_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_29_io_in_weight = PE_Array_23_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_29_io_in_psum = PE_Array_23_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_30_clock = clock;
  assign PE_Array_24_30_reset = reset;
  assign PE_Array_24_30_io_in_activate = PE_Array_24_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_30_io_in_weight = PE_Array_23_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_30_io_in_psum = PE_Array_23_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_24_31_clock = clock;
  assign PE_Array_24_31_reset = reset;
  assign PE_Array_24_31_io_in_activate = PE_Array_24_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_24_31_io_in_weight = PE_Array_23_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_24_31_io_in_psum = PE_Array_23_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_24_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_24_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_0_clock = clock;
  assign PE_Array_25_0_reset = reset;
  assign PE_Array_25_0_io_in_activate = io_activate_25; // @[DataPath.scala 11:26]
  assign PE_Array_25_0_io_in_weight = PE_Array_24_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_0_io_in_psum = PE_Array_24_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_1_clock = clock;
  assign PE_Array_25_1_reset = reset;
  assign PE_Array_25_1_io_in_activate = PE_Array_25_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_1_io_in_weight = PE_Array_24_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_1_io_in_psum = PE_Array_24_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_2_clock = clock;
  assign PE_Array_25_2_reset = reset;
  assign PE_Array_25_2_io_in_activate = PE_Array_25_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_2_io_in_weight = PE_Array_24_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_2_io_in_psum = PE_Array_24_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_3_clock = clock;
  assign PE_Array_25_3_reset = reset;
  assign PE_Array_25_3_io_in_activate = PE_Array_25_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_3_io_in_weight = PE_Array_24_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_3_io_in_psum = PE_Array_24_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_4_clock = clock;
  assign PE_Array_25_4_reset = reset;
  assign PE_Array_25_4_io_in_activate = PE_Array_25_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_4_io_in_weight = PE_Array_24_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_4_io_in_psum = PE_Array_24_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_5_clock = clock;
  assign PE_Array_25_5_reset = reset;
  assign PE_Array_25_5_io_in_activate = PE_Array_25_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_5_io_in_weight = PE_Array_24_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_5_io_in_psum = PE_Array_24_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_6_clock = clock;
  assign PE_Array_25_6_reset = reset;
  assign PE_Array_25_6_io_in_activate = PE_Array_25_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_6_io_in_weight = PE_Array_24_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_6_io_in_psum = PE_Array_24_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_7_clock = clock;
  assign PE_Array_25_7_reset = reset;
  assign PE_Array_25_7_io_in_activate = PE_Array_25_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_7_io_in_weight = PE_Array_24_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_7_io_in_psum = PE_Array_24_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_8_clock = clock;
  assign PE_Array_25_8_reset = reset;
  assign PE_Array_25_8_io_in_activate = PE_Array_25_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_8_io_in_weight = PE_Array_24_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_8_io_in_psum = PE_Array_24_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_9_clock = clock;
  assign PE_Array_25_9_reset = reset;
  assign PE_Array_25_9_io_in_activate = PE_Array_25_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_9_io_in_weight = PE_Array_24_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_9_io_in_psum = PE_Array_24_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_10_clock = clock;
  assign PE_Array_25_10_reset = reset;
  assign PE_Array_25_10_io_in_activate = PE_Array_25_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_10_io_in_weight = PE_Array_24_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_10_io_in_psum = PE_Array_24_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_11_clock = clock;
  assign PE_Array_25_11_reset = reset;
  assign PE_Array_25_11_io_in_activate = PE_Array_25_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_11_io_in_weight = PE_Array_24_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_11_io_in_psum = PE_Array_24_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_12_clock = clock;
  assign PE_Array_25_12_reset = reset;
  assign PE_Array_25_12_io_in_activate = PE_Array_25_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_12_io_in_weight = PE_Array_24_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_12_io_in_psum = PE_Array_24_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_13_clock = clock;
  assign PE_Array_25_13_reset = reset;
  assign PE_Array_25_13_io_in_activate = PE_Array_25_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_13_io_in_weight = PE_Array_24_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_13_io_in_psum = PE_Array_24_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_14_clock = clock;
  assign PE_Array_25_14_reset = reset;
  assign PE_Array_25_14_io_in_activate = PE_Array_25_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_14_io_in_weight = PE_Array_24_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_14_io_in_psum = PE_Array_24_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_15_clock = clock;
  assign PE_Array_25_15_reset = reset;
  assign PE_Array_25_15_io_in_activate = PE_Array_25_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_15_io_in_weight = PE_Array_24_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_15_io_in_psum = PE_Array_24_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_16_clock = clock;
  assign PE_Array_25_16_reset = reset;
  assign PE_Array_25_16_io_in_activate = PE_Array_25_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_16_io_in_weight = PE_Array_24_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_16_io_in_psum = PE_Array_24_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_17_clock = clock;
  assign PE_Array_25_17_reset = reset;
  assign PE_Array_25_17_io_in_activate = PE_Array_25_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_17_io_in_weight = PE_Array_24_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_17_io_in_psum = PE_Array_24_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_18_clock = clock;
  assign PE_Array_25_18_reset = reset;
  assign PE_Array_25_18_io_in_activate = PE_Array_25_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_18_io_in_weight = PE_Array_24_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_18_io_in_psum = PE_Array_24_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_19_clock = clock;
  assign PE_Array_25_19_reset = reset;
  assign PE_Array_25_19_io_in_activate = PE_Array_25_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_19_io_in_weight = PE_Array_24_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_19_io_in_psum = PE_Array_24_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_20_clock = clock;
  assign PE_Array_25_20_reset = reset;
  assign PE_Array_25_20_io_in_activate = PE_Array_25_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_20_io_in_weight = PE_Array_24_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_20_io_in_psum = PE_Array_24_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_21_clock = clock;
  assign PE_Array_25_21_reset = reset;
  assign PE_Array_25_21_io_in_activate = PE_Array_25_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_21_io_in_weight = PE_Array_24_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_21_io_in_psum = PE_Array_24_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_22_clock = clock;
  assign PE_Array_25_22_reset = reset;
  assign PE_Array_25_22_io_in_activate = PE_Array_25_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_22_io_in_weight = PE_Array_24_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_22_io_in_psum = PE_Array_24_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_23_clock = clock;
  assign PE_Array_25_23_reset = reset;
  assign PE_Array_25_23_io_in_activate = PE_Array_25_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_23_io_in_weight = PE_Array_24_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_23_io_in_psum = PE_Array_24_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_24_clock = clock;
  assign PE_Array_25_24_reset = reset;
  assign PE_Array_25_24_io_in_activate = PE_Array_25_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_24_io_in_weight = PE_Array_24_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_24_io_in_psum = PE_Array_24_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_25_clock = clock;
  assign PE_Array_25_25_reset = reset;
  assign PE_Array_25_25_io_in_activate = PE_Array_25_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_25_io_in_weight = PE_Array_24_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_25_io_in_psum = PE_Array_24_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_26_clock = clock;
  assign PE_Array_25_26_reset = reset;
  assign PE_Array_25_26_io_in_activate = PE_Array_25_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_26_io_in_weight = PE_Array_24_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_26_io_in_psum = PE_Array_24_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_27_clock = clock;
  assign PE_Array_25_27_reset = reset;
  assign PE_Array_25_27_io_in_activate = PE_Array_25_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_27_io_in_weight = PE_Array_24_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_27_io_in_psum = PE_Array_24_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_28_clock = clock;
  assign PE_Array_25_28_reset = reset;
  assign PE_Array_25_28_io_in_activate = PE_Array_25_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_28_io_in_weight = PE_Array_24_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_28_io_in_psum = PE_Array_24_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_29_clock = clock;
  assign PE_Array_25_29_reset = reset;
  assign PE_Array_25_29_io_in_activate = PE_Array_25_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_29_io_in_weight = PE_Array_24_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_29_io_in_psum = PE_Array_24_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_30_clock = clock;
  assign PE_Array_25_30_reset = reset;
  assign PE_Array_25_30_io_in_activate = PE_Array_25_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_30_io_in_weight = PE_Array_24_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_30_io_in_psum = PE_Array_24_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_25_31_clock = clock;
  assign PE_Array_25_31_reset = reset;
  assign PE_Array_25_31_io_in_activate = PE_Array_25_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_25_31_io_in_weight = PE_Array_24_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_25_31_io_in_psum = PE_Array_24_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_25_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_25_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_0_clock = clock;
  assign PE_Array_26_0_reset = reset;
  assign PE_Array_26_0_io_in_activate = io_activate_26; // @[DataPath.scala 11:26]
  assign PE_Array_26_0_io_in_weight = PE_Array_25_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_0_io_in_psum = PE_Array_25_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_1_clock = clock;
  assign PE_Array_26_1_reset = reset;
  assign PE_Array_26_1_io_in_activate = PE_Array_26_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_1_io_in_weight = PE_Array_25_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_1_io_in_psum = PE_Array_25_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_2_clock = clock;
  assign PE_Array_26_2_reset = reset;
  assign PE_Array_26_2_io_in_activate = PE_Array_26_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_2_io_in_weight = PE_Array_25_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_2_io_in_psum = PE_Array_25_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_3_clock = clock;
  assign PE_Array_26_3_reset = reset;
  assign PE_Array_26_3_io_in_activate = PE_Array_26_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_3_io_in_weight = PE_Array_25_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_3_io_in_psum = PE_Array_25_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_4_clock = clock;
  assign PE_Array_26_4_reset = reset;
  assign PE_Array_26_4_io_in_activate = PE_Array_26_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_4_io_in_weight = PE_Array_25_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_4_io_in_psum = PE_Array_25_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_5_clock = clock;
  assign PE_Array_26_5_reset = reset;
  assign PE_Array_26_5_io_in_activate = PE_Array_26_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_5_io_in_weight = PE_Array_25_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_5_io_in_psum = PE_Array_25_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_6_clock = clock;
  assign PE_Array_26_6_reset = reset;
  assign PE_Array_26_6_io_in_activate = PE_Array_26_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_6_io_in_weight = PE_Array_25_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_6_io_in_psum = PE_Array_25_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_7_clock = clock;
  assign PE_Array_26_7_reset = reset;
  assign PE_Array_26_7_io_in_activate = PE_Array_26_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_7_io_in_weight = PE_Array_25_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_7_io_in_psum = PE_Array_25_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_8_clock = clock;
  assign PE_Array_26_8_reset = reset;
  assign PE_Array_26_8_io_in_activate = PE_Array_26_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_8_io_in_weight = PE_Array_25_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_8_io_in_psum = PE_Array_25_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_9_clock = clock;
  assign PE_Array_26_9_reset = reset;
  assign PE_Array_26_9_io_in_activate = PE_Array_26_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_9_io_in_weight = PE_Array_25_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_9_io_in_psum = PE_Array_25_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_10_clock = clock;
  assign PE_Array_26_10_reset = reset;
  assign PE_Array_26_10_io_in_activate = PE_Array_26_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_10_io_in_weight = PE_Array_25_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_10_io_in_psum = PE_Array_25_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_11_clock = clock;
  assign PE_Array_26_11_reset = reset;
  assign PE_Array_26_11_io_in_activate = PE_Array_26_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_11_io_in_weight = PE_Array_25_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_11_io_in_psum = PE_Array_25_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_12_clock = clock;
  assign PE_Array_26_12_reset = reset;
  assign PE_Array_26_12_io_in_activate = PE_Array_26_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_12_io_in_weight = PE_Array_25_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_12_io_in_psum = PE_Array_25_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_13_clock = clock;
  assign PE_Array_26_13_reset = reset;
  assign PE_Array_26_13_io_in_activate = PE_Array_26_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_13_io_in_weight = PE_Array_25_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_13_io_in_psum = PE_Array_25_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_14_clock = clock;
  assign PE_Array_26_14_reset = reset;
  assign PE_Array_26_14_io_in_activate = PE_Array_26_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_14_io_in_weight = PE_Array_25_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_14_io_in_psum = PE_Array_25_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_15_clock = clock;
  assign PE_Array_26_15_reset = reset;
  assign PE_Array_26_15_io_in_activate = PE_Array_26_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_15_io_in_weight = PE_Array_25_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_15_io_in_psum = PE_Array_25_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_16_clock = clock;
  assign PE_Array_26_16_reset = reset;
  assign PE_Array_26_16_io_in_activate = PE_Array_26_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_16_io_in_weight = PE_Array_25_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_16_io_in_psum = PE_Array_25_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_17_clock = clock;
  assign PE_Array_26_17_reset = reset;
  assign PE_Array_26_17_io_in_activate = PE_Array_26_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_17_io_in_weight = PE_Array_25_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_17_io_in_psum = PE_Array_25_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_18_clock = clock;
  assign PE_Array_26_18_reset = reset;
  assign PE_Array_26_18_io_in_activate = PE_Array_26_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_18_io_in_weight = PE_Array_25_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_18_io_in_psum = PE_Array_25_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_19_clock = clock;
  assign PE_Array_26_19_reset = reset;
  assign PE_Array_26_19_io_in_activate = PE_Array_26_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_19_io_in_weight = PE_Array_25_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_19_io_in_psum = PE_Array_25_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_20_clock = clock;
  assign PE_Array_26_20_reset = reset;
  assign PE_Array_26_20_io_in_activate = PE_Array_26_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_20_io_in_weight = PE_Array_25_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_20_io_in_psum = PE_Array_25_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_21_clock = clock;
  assign PE_Array_26_21_reset = reset;
  assign PE_Array_26_21_io_in_activate = PE_Array_26_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_21_io_in_weight = PE_Array_25_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_21_io_in_psum = PE_Array_25_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_22_clock = clock;
  assign PE_Array_26_22_reset = reset;
  assign PE_Array_26_22_io_in_activate = PE_Array_26_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_22_io_in_weight = PE_Array_25_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_22_io_in_psum = PE_Array_25_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_23_clock = clock;
  assign PE_Array_26_23_reset = reset;
  assign PE_Array_26_23_io_in_activate = PE_Array_26_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_23_io_in_weight = PE_Array_25_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_23_io_in_psum = PE_Array_25_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_24_clock = clock;
  assign PE_Array_26_24_reset = reset;
  assign PE_Array_26_24_io_in_activate = PE_Array_26_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_24_io_in_weight = PE_Array_25_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_24_io_in_psum = PE_Array_25_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_25_clock = clock;
  assign PE_Array_26_25_reset = reset;
  assign PE_Array_26_25_io_in_activate = PE_Array_26_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_25_io_in_weight = PE_Array_25_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_25_io_in_psum = PE_Array_25_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_26_clock = clock;
  assign PE_Array_26_26_reset = reset;
  assign PE_Array_26_26_io_in_activate = PE_Array_26_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_26_io_in_weight = PE_Array_25_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_26_io_in_psum = PE_Array_25_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_27_clock = clock;
  assign PE_Array_26_27_reset = reset;
  assign PE_Array_26_27_io_in_activate = PE_Array_26_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_27_io_in_weight = PE_Array_25_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_27_io_in_psum = PE_Array_25_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_28_clock = clock;
  assign PE_Array_26_28_reset = reset;
  assign PE_Array_26_28_io_in_activate = PE_Array_26_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_28_io_in_weight = PE_Array_25_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_28_io_in_psum = PE_Array_25_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_29_clock = clock;
  assign PE_Array_26_29_reset = reset;
  assign PE_Array_26_29_io_in_activate = PE_Array_26_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_29_io_in_weight = PE_Array_25_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_29_io_in_psum = PE_Array_25_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_30_clock = clock;
  assign PE_Array_26_30_reset = reset;
  assign PE_Array_26_30_io_in_activate = PE_Array_26_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_30_io_in_weight = PE_Array_25_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_30_io_in_psum = PE_Array_25_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_26_31_clock = clock;
  assign PE_Array_26_31_reset = reset;
  assign PE_Array_26_31_io_in_activate = PE_Array_26_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_26_31_io_in_weight = PE_Array_25_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_26_31_io_in_psum = PE_Array_25_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_26_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_26_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_0_clock = clock;
  assign PE_Array_27_0_reset = reset;
  assign PE_Array_27_0_io_in_activate = io_activate_27; // @[DataPath.scala 11:26]
  assign PE_Array_27_0_io_in_weight = PE_Array_26_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_0_io_in_psum = PE_Array_26_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_1_clock = clock;
  assign PE_Array_27_1_reset = reset;
  assign PE_Array_27_1_io_in_activate = PE_Array_27_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_1_io_in_weight = PE_Array_26_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_1_io_in_psum = PE_Array_26_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_2_clock = clock;
  assign PE_Array_27_2_reset = reset;
  assign PE_Array_27_2_io_in_activate = PE_Array_27_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_2_io_in_weight = PE_Array_26_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_2_io_in_psum = PE_Array_26_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_3_clock = clock;
  assign PE_Array_27_3_reset = reset;
  assign PE_Array_27_3_io_in_activate = PE_Array_27_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_3_io_in_weight = PE_Array_26_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_3_io_in_psum = PE_Array_26_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_4_clock = clock;
  assign PE_Array_27_4_reset = reset;
  assign PE_Array_27_4_io_in_activate = PE_Array_27_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_4_io_in_weight = PE_Array_26_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_4_io_in_psum = PE_Array_26_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_5_clock = clock;
  assign PE_Array_27_5_reset = reset;
  assign PE_Array_27_5_io_in_activate = PE_Array_27_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_5_io_in_weight = PE_Array_26_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_5_io_in_psum = PE_Array_26_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_6_clock = clock;
  assign PE_Array_27_6_reset = reset;
  assign PE_Array_27_6_io_in_activate = PE_Array_27_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_6_io_in_weight = PE_Array_26_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_6_io_in_psum = PE_Array_26_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_7_clock = clock;
  assign PE_Array_27_7_reset = reset;
  assign PE_Array_27_7_io_in_activate = PE_Array_27_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_7_io_in_weight = PE_Array_26_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_7_io_in_psum = PE_Array_26_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_8_clock = clock;
  assign PE_Array_27_8_reset = reset;
  assign PE_Array_27_8_io_in_activate = PE_Array_27_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_8_io_in_weight = PE_Array_26_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_8_io_in_psum = PE_Array_26_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_9_clock = clock;
  assign PE_Array_27_9_reset = reset;
  assign PE_Array_27_9_io_in_activate = PE_Array_27_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_9_io_in_weight = PE_Array_26_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_9_io_in_psum = PE_Array_26_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_10_clock = clock;
  assign PE_Array_27_10_reset = reset;
  assign PE_Array_27_10_io_in_activate = PE_Array_27_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_10_io_in_weight = PE_Array_26_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_10_io_in_psum = PE_Array_26_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_11_clock = clock;
  assign PE_Array_27_11_reset = reset;
  assign PE_Array_27_11_io_in_activate = PE_Array_27_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_11_io_in_weight = PE_Array_26_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_11_io_in_psum = PE_Array_26_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_12_clock = clock;
  assign PE_Array_27_12_reset = reset;
  assign PE_Array_27_12_io_in_activate = PE_Array_27_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_12_io_in_weight = PE_Array_26_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_12_io_in_psum = PE_Array_26_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_13_clock = clock;
  assign PE_Array_27_13_reset = reset;
  assign PE_Array_27_13_io_in_activate = PE_Array_27_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_13_io_in_weight = PE_Array_26_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_13_io_in_psum = PE_Array_26_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_14_clock = clock;
  assign PE_Array_27_14_reset = reset;
  assign PE_Array_27_14_io_in_activate = PE_Array_27_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_14_io_in_weight = PE_Array_26_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_14_io_in_psum = PE_Array_26_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_15_clock = clock;
  assign PE_Array_27_15_reset = reset;
  assign PE_Array_27_15_io_in_activate = PE_Array_27_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_15_io_in_weight = PE_Array_26_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_15_io_in_psum = PE_Array_26_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_16_clock = clock;
  assign PE_Array_27_16_reset = reset;
  assign PE_Array_27_16_io_in_activate = PE_Array_27_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_16_io_in_weight = PE_Array_26_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_16_io_in_psum = PE_Array_26_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_17_clock = clock;
  assign PE_Array_27_17_reset = reset;
  assign PE_Array_27_17_io_in_activate = PE_Array_27_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_17_io_in_weight = PE_Array_26_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_17_io_in_psum = PE_Array_26_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_18_clock = clock;
  assign PE_Array_27_18_reset = reset;
  assign PE_Array_27_18_io_in_activate = PE_Array_27_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_18_io_in_weight = PE_Array_26_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_18_io_in_psum = PE_Array_26_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_19_clock = clock;
  assign PE_Array_27_19_reset = reset;
  assign PE_Array_27_19_io_in_activate = PE_Array_27_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_19_io_in_weight = PE_Array_26_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_19_io_in_psum = PE_Array_26_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_20_clock = clock;
  assign PE_Array_27_20_reset = reset;
  assign PE_Array_27_20_io_in_activate = PE_Array_27_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_20_io_in_weight = PE_Array_26_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_20_io_in_psum = PE_Array_26_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_21_clock = clock;
  assign PE_Array_27_21_reset = reset;
  assign PE_Array_27_21_io_in_activate = PE_Array_27_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_21_io_in_weight = PE_Array_26_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_21_io_in_psum = PE_Array_26_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_22_clock = clock;
  assign PE_Array_27_22_reset = reset;
  assign PE_Array_27_22_io_in_activate = PE_Array_27_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_22_io_in_weight = PE_Array_26_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_22_io_in_psum = PE_Array_26_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_23_clock = clock;
  assign PE_Array_27_23_reset = reset;
  assign PE_Array_27_23_io_in_activate = PE_Array_27_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_23_io_in_weight = PE_Array_26_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_23_io_in_psum = PE_Array_26_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_24_clock = clock;
  assign PE_Array_27_24_reset = reset;
  assign PE_Array_27_24_io_in_activate = PE_Array_27_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_24_io_in_weight = PE_Array_26_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_24_io_in_psum = PE_Array_26_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_25_clock = clock;
  assign PE_Array_27_25_reset = reset;
  assign PE_Array_27_25_io_in_activate = PE_Array_27_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_25_io_in_weight = PE_Array_26_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_25_io_in_psum = PE_Array_26_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_26_clock = clock;
  assign PE_Array_27_26_reset = reset;
  assign PE_Array_27_26_io_in_activate = PE_Array_27_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_26_io_in_weight = PE_Array_26_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_26_io_in_psum = PE_Array_26_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_27_clock = clock;
  assign PE_Array_27_27_reset = reset;
  assign PE_Array_27_27_io_in_activate = PE_Array_27_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_27_io_in_weight = PE_Array_26_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_27_io_in_psum = PE_Array_26_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_28_clock = clock;
  assign PE_Array_27_28_reset = reset;
  assign PE_Array_27_28_io_in_activate = PE_Array_27_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_28_io_in_weight = PE_Array_26_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_28_io_in_psum = PE_Array_26_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_29_clock = clock;
  assign PE_Array_27_29_reset = reset;
  assign PE_Array_27_29_io_in_activate = PE_Array_27_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_29_io_in_weight = PE_Array_26_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_29_io_in_psum = PE_Array_26_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_30_clock = clock;
  assign PE_Array_27_30_reset = reset;
  assign PE_Array_27_30_io_in_activate = PE_Array_27_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_30_io_in_weight = PE_Array_26_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_30_io_in_psum = PE_Array_26_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_27_31_clock = clock;
  assign PE_Array_27_31_reset = reset;
  assign PE_Array_27_31_io_in_activate = PE_Array_27_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_27_31_io_in_weight = PE_Array_26_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_27_31_io_in_psum = PE_Array_26_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_27_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_27_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_0_clock = clock;
  assign PE_Array_28_0_reset = reset;
  assign PE_Array_28_0_io_in_activate = io_activate_28; // @[DataPath.scala 11:26]
  assign PE_Array_28_0_io_in_weight = PE_Array_27_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_0_io_in_psum = PE_Array_27_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_1_clock = clock;
  assign PE_Array_28_1_reset = reset;
  assign PE_Array_28_1_io_in_activate = PE_Array_28_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_1_io_in_weight = PE_Array_27_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_1_io_in_psum = PE_Array_27_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_2_clock = clock;
  assign PE_Array_28_2_reset = reset;
  assign PE_Array_28_2_io_in_activate = PE_Array_28_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_2_io_in_weight = PE_Array_27_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_2_io_in_psum = PE_Array_27_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_3_clock = clock;
  assign PE_Array_28_3_reset = reset;
  assign PE_Array_28_3_io_in_activate = PE_Array_28_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_3_io_in_weight = PE_Array_27_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_3_io_in_psum = PE_Array_27_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_4_clock = clock;
  assign PE_Array_28_4_reset = reset;
  assign PE_Array_28_4_io_in_activate = PE_Array_28_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_4_io_in_weight = PE_Array_27_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_4_io_in_psum = PE_Array_27_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_5_clock = clock;
  assign PE_Array_28_5_reset = reset;
  assign PE_Array_28_5_io_in_activate = PE_Array_28_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_5_io_in_weight = PE_Array_27_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_5_io_in_psum = PE_Array_27_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_6_clock = clock;
  assign PE_Array_28_6_reset = reset;
  assign PE_Array_28_6_io_in_activate = PE_Array_28_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_6_io_in_weight = PE_Array_27_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_6_io_in_psum = PE_Array_27_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_7_clock = clock;
  assign PE_Array_28_7_reset = reset;
  assign PE_Array_28_7_io_in_activate = PE_Array_28_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_7_io_in_weight = PE_Array_27_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_7_io_in_psum = PE_Array_27_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_8_clock = clock;
  assign PE_Array_28_8_reset = reset;
  assign PE_Array_28_8_io_in_activate = PE_Array_28_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_8_io_in_weight = PE_Array_27_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_8_io_in_psum = PE_Array_27_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_9_clock = clock;
  assign PE_Array_28_9_reset = reset;
  assign PE_Array_28_9_io_in_activate = PE_Array_28_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_9_io_in_weight = PE_Array_27_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_9_io_in_psum = PE_Array_27_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_10_clock = clock;
  assign PE_Array_28_10_reset = reset;
  assign PE_Array_28_10_io_in_activate = PE_Array_28_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_10_io_in_weight = PE_Array_27_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_10_io_in_psum = PE_Array_27_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_11_clock = clock;
  assign PE_Array_28_11_reset = reset;
  assign PE_Array_28_11_io_in_activate = PE_Array_28_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_11_io_in_weight = PE_Array_27_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_11_io_in_psum = PE_Array_27_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_12_clock = clock;
  assign PE_Array_28_12_reset = reset;
  assign PE_Array_28_12_io_in_activate = PE_Array_28_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_12_io_in_weight = PE_Array_27_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_12_io_in_psum = PE_Array_27_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_13_clock = clock;
  assign PE_Array_28_13_reset = reset;
  assign PE_Array_28_13_io_in_activate = PE_Array_28_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_13_io_in_weight = PE_Array_27_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_13_io_in_psum = PE_Array_27_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_14_clock = clock;
  assign PE_Array_28_14_reset = reset;
  assign PE_Array_28_14_io_in_activate = PE_Array_28_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_14_io_in_weight = PE_Array_27_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_14_io_in_psum = PE_Array_27_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_15_clock = clock;
  assign PE_Array_28_15_reset = reset;
  assign PE_Array_28_15_io_in_activate = PE_Array_28_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_15_io_in_weight = PE_Array_27_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_15_io_in_psum = PE_Array_27_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_16_clock = clock;
  assign PE_Array_28_16_reset = reset;
  assign PE_Array_28_16_io_in_activate = PE_Array_28_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_16_io_in_weight = PE_Array_27_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_16_io_in_psum = PE_Array_27_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_17_clock = clock;
  assign PE_Array_28_17_reset = reset;
  assign PE_Array_28_17_io_in_activate = PE_Array_28_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_17_io_in_weight = PE_Array_27_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_17_io_in_psum = PE_Array_27_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_18_clock = clock;
  assign PE_Array_28_18_reset = reset;
  assign PE_Array_28_18_io_in_activate = PE_Array_28_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_18_io_in_weight = PE_Array_27_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_18_io_in_psum = PE_Array_27_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_19_clock = clock;
  assign PE_Array_28_19_reset = reset;
  assign PE_Array_28_19_io_in_activate = PE_Array_28_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_19_io_in_weight = PE_Array_27_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_19_io_in_psum = PE_Array_27_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_20_clock = clock;
  assign PE_Array_28_20_reset = reset;
  assign PE_Array_28_20_io_in_activate = PE_Array_28_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_20_io_in_weight = PE_Array_27_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_20_io_in_psum = PE_Array_27_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_21_clock = clock;
  assign PE_Array_28_21_reset = reset;
  assign PE_Array_28_21_io_in_activate = PE_Array_28_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_21_io_in_weight = PE_Array_27_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_21_io_in_psum = PE_Array_27_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_22_clock = clock;
  assign PE_Array_28_22_reset = reset;
  assign PE_Array_28_22_io_in_activate = PE_Array_28_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_22_io_in_weight = PE_Array_27_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_22_io_in_psum = PE_Array_27_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_23_clock = clock;
  assign PE_Array_28_23_reset = reset;
  assign PE_Array_28_23_io_in_activate = PE_Array_28_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_23_io_in_weight = PE_Array_27_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_23_io_in_psum = PE_Array_27_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_24_clock = clock;
  assign PE_Array_28_24_reset = reset;
  assign PE_Array_28_24_io_in_activate = PE_Array_28_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_24_io_in_weight = PE_Array_27_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_24_io_in_psum = PE_Array_27_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_25_clock = clock;
  assign PE_Array_28_25_reset = reset;
  assign PE_Array_28_25_io_in_activate = PE_Array_28_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_25_io_in_weight = PE_Array_27_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_25_io_in_psum = PE_Array_27_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_26_clock = clock;
  assign PE_Array_28_26_reset = reset;
  assign PE_Array_28_26_io_in_activate = PE_Array_28_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_26_io_in_weight = PE_Array_27_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_26_io_in_psum = PE_Array_27_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_27_clock = clock;
  assign PE_Array_28_27_reset = reset;
  assign PE_Array_28_27_io_in_activate = PE_Array_28_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_27_io_in_weight = PE_Array_27_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_27_io_in_psum = PE_Array_27_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_28_clock = clock;
  assign PE_Array_28_28_reset = reset;
  assign PE_Array_28_28_io_in_activate = PE_Array_28_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_28_io_in_weight = PE_Array_27_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_28_io_in_psum = PE_Array_27_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_29_clock = clock;
  assign PE_Array_28_29_reset = reset;
  assign PE_Array_28_29_io_in_activate = PE_Array_28_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_29_io_in_weight = PE_Array_27_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_29_io_in_psum = PE_Array_27_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_30_clock = clock;
  assign PE_Array_28_30_reset = reset;
  assign PE_Array_28_30_io_in_activate = PE_Array_28_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_30_io_in_weight = PE_Array_27_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_30_io_in_psum = PE_Array_27_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_28_31_clock = clock;
  assign PE_Array_28_31_reset = reset;
  assign PE_Array_28_31_io_in_activate = PE_Array_28_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_28_31_io_in_weight = PE_Array_27_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_28_31_io_in_psum = PE_Array_27_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_28_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_28_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_0_clock = clock;
  assign PE_Array_29_0_reset = reset;
  assign PE_Array_29_0_io_in_activate = io_activate_29; // @[DataPath.scala 11:26]
  assign PE_Array_29_0_io_in_weight = PE_Array_28_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_0_io_in_psum = PE_Array_28_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_1_clock = clock;
  assign PE_Array_29_1_reset = reset;
  assign PE_Array_29_1_io_in_activate = PE_Array_29_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_1_io_in_weight = PE_Array_28_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_1_io_in_psum = PE_Array_28_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_2_clock = clock;
  assign PE_Array_29_2_reset = reset;
  assign PE_Array_29_2_io_in_activate = PE_Array_29_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_2_io_in_weight = PE_Array_28_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_2_io_in_psum = PE_Array_28_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_3_clock = clock;
  assign PE_Array_29_3_reset = reset;
  assign PE_Array_29_3_io_in_activate = PE_Array_29_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_3_io_in_weight = PE_Array_28_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_3_io_in_psum = PE_Array_28_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_4_clock = clock;
  assign PE_Array_29_4_reset = reset;
  assign PE_Array_29_4_io_in_activate = PE_Array_29_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_4_io_in_weight = PE_Array_28_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_4_io_in_psum = PE_Array_28_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_5_clock = clock;
  assign PE_Array_29_5_reset = reset;
  assign PE_Array_29_5_io_in_activate = PE_Array_29_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_5_io_in_weight = PE_Array_28_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_5_io_in_psum = PE_Array_28_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_6_clock = clock;
  assign PE_Array_29_6_reset = reset;
  assign PE_Array_29_6_io_in_activate = PE_Array_29_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_6_io_in_weight = PE_Array_28_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_6_io_in_psum = PE_Array_28_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_7_clock = clock;
  assign PE_Array_29_7_reset = reset;
  assign PE_Array_29_7_io_in_activate = PE_Array_29_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_7_io_in_weight = PE_Array_28_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_7_io_in_psum = PE_Array_28_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_8_clock = clock;
  assign PE_Array_29_8_reset = reset;
  assign PE_Array_29_8_io_in_activate = PE_Array_29_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_8_io_in_weight = PE_Array_28_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_8_io_in_psum = PE_Array_28_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_9_clock = clock;
  assign PE_Array_29_9_reset = reset;
  assign PE_Array_29_9_io_in_activate = PE_Array_29_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_9_io_in_weight = PE_Array_28_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_9_io_in_psum = PE_Array_28_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_10_clock = clock;
  assign PE_Array_29_10_reset = reset;
  assign PE_Array_29_10_io_in_activate = PE_Array_29_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_10_io_in_weight = PE_Array_28_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_10_io_in_psum = PE_Array_28_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_11_clock = clock;
  assign PE_Array_29_11_reset = reset;
  assign PE_Array_29_11_io_in_activate = PE_Array_29_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_11_io_in_weight = PE_Array_28_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_11_io_in_psum = PE_Array_28_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_12_clock = clock;
  assign PE_Array_29_12_reset = reset;
  assign PE_Array_29_12_io_in_activate = PE_Array_29_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_12_io_in_weight = PE_Array_28_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_12_io_in_psum = PE_Array_28_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_13_clock = clock;
  assign PE_Array_29_13_reset = reset;
  assign PE_Array_29_13_io_in_activate = PE_Array_29_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_13_io_in_weight = PE_Array_28_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_13_io_in_psum = PE_Array_28_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_14_clock = clock;
  assign PE_Array_29_14_reset = reset;
  assign PE_Array_29_14_io_in_activate = PE_Array_29_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_14_io_in_weight = PE_Array_28_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_14_io_in_psum = PE_Array_28_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_15_clock = clock;
  assign PE_Array_29_15_reset = reset;
  assign PE_Array_29_15_io_in_activate = PE_Array_29_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_15_io_in_weight = PE_Array_28_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_15_io_in_psum = PE_Array_28_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_16_clock = clock;
  assign PE_Array_29_16_reset = reset;
  assign PE_Array_29_16_io_in_activate = PE_Array_29_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_16_io_in_weight = PE_Array_28_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_16_io_in_psum = PE_Array_28_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_17_clock = clock;
  assign PE_Array_29_17_reset = reset;
  assign PE_Array_29_17_io_in_activate = PE_Array_29_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_17_io_in_weight = PE_Array_28_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_17_io_in_psum = PE_Array_28_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_18_clock = clock;
  assign PE_Array_29_18_reset = reset;
  assign PE_Array_29_18_io_in_activate = PE_Array_29_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_18_io_in_weight = PE_Array_28_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_18_io_in_psum = PE_Array_28_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_19_clock = clock;
  assign PE_Array_29_19_reset = reset;
  assign PE_Array_29_19_io_in_activate = PE_Array_29_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_19_io_in_weight = PE_Array_28_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_19_io_in_psum = PE_Array_28_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_20_clock = clock;
  assign PE_Array_29_20_reset = reset;
  assign PE_Array_29_20_io_in_activate = PE_Array_29_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_20_io_in_weight = PE_Array_28_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_20_io_in_psum = PE_Array_28_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_21_clock = clock;
  assign PE_Array_29_21_reset = reset;
  assign PE_Array_29_21_io_in_activate = PE_Array_29_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_21_io_in_weight = PE_Array_28_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_21_io_in_psum = PE_Array_28_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_22_clock = clock;
  assign PE_Array_29_22_reset = reset;
  assign PE_Array_29_22_io_in_activate = PE_Array_29_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_22_io_in_weight = PE_Array_28_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_22_io_in_psum = PE_Array_28_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_23_clock = clock;
  assign PE_Array_29_23_reset = reset;
  assign PE_Array_29_23_io_in_activate = PE_Array_29_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_23_io_in_weight = PE_Array_28_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_23_io_in_psum = PE_Array_28_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_24_clock = clock;
  assign PE_Array_29_24_reset = reset;
  assign PE_Array_29_24_io_in_activate = PE_Array_29_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_24_io_in_weight = PE_Array_28_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_24_io_in_psum = PE_Array_28_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_25_clock = clock;
  assign PE_Array_29_25_reset = reset;
  assign PE_Array_29_25_io_in_activate = PE_Array_29_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_25_io_in_weight = PE_Array_28_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_25_io_in_psum = PE_Array_28_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_26_clock = clock;
  assign PE_Array_29_26_reset = reset;
  assign PE_Array_29_26_io_in_activate = PE_Array_29_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_26_io_in_weight = PE_Array_28_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_26_io_in_psum = PE_Array_28_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_27_clock = clock;
  assign PE_Array_29_27_reset = reset;
  assign PE_Array_29_27_io_in_activate = PE_Array_29_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_27_io_in_weight = PE_Array_28_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_27_io_in_psum = PE_Array_28_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_28_clock = clock;
  assign PE_Array_29_28_reset = reset;
  assign PE_Array_29_28_io_in_activate = PE_Array_29_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_28_io_in_weight = PE_Array_28_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_28_io_in_psum = PE_Array_28_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_29_clock = clock;
  assign PE_Array_29_29_reset = reset;
  assign PE_Array_29_29_io_in_activate = PE_Array_29_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_29_io_in_weight = PE_Array_28_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_29_io_in_psum = PE_Array_28_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_30_clock = clock;
  assign PE_Array_29_30_reset = reset;
  assign PE_Array_29_30_io_in_activate = PE_Array_29_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_30_io_in_weight = PE_Array_28_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_30_io_in_psum = PE_Array_28_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_29_31_clock = clock;
  assign PE_Array_29_31_reset = reset;
  assign PE_Array_29_31_io_in_activate = PE_Array_29_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_29_31_io_in_weight = PE_Array_28_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_29_31_io_in_psum = PE_Array_28_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_29_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_29_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_0_clock = clock;
  assign PE_Array_30_0_reset = reset;
  assign PE_Array_30_0_io_in_activate = io_activate_30; // @[DataPath.scala 11:26]
  assign PE_Array_30_0_io_in_weight = PE_Array_29_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_0_io_in_psum = PE_Array_29_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_1_clock = clock;
  assign PE_Array_30_1_reset = reset;
  assign PE_Array_30_1_io_in_activate = PE_Array_30_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_1_io_in_weight = PE_Array_29_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_1_io_in_psum = PE_Array_29_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_2_clock = clock;
  assign PE_Array_30_2_reset = reset;
  assign PE_Array_30_2_io_in_activate = PE_Array_30_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_2_io_in_weight = PE_Array_29_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_2_io_in_psum = PE_Array_29_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_3_clock = clock;
  assign PE_Array_30_3_reset = reset;
  assign PE_Array_30_3_io_in_activate = PE_Array_30_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_3_io_in_weight = PE_Array_29_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_3_io_in_psum = PE_Array_29_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_4_clock = clock;
  assign PE_Array_30_4_reset = reset;
  assign PE_Array_30_4_io_in_activate = PE_Array_30_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_4_io_in_weight = PE_Array_29_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_4_io_in_psum = PE_Array_29_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_5_clock = clock;
  assign PE_Array_30_5_reset = reset;
  assign PE_Array_30_5_io_in_activate = PE_Array_30_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_5_io_in_weight = PE_Array_29_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_5_io_in_psum = PE_Array_29_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_6_clock = clock;
  assign PE_Array_30_6_reset = reset;
  assign PE_Array_30_6_io_in_activate = PE_Array_30_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_6_io_in_weight = PE_Array_29_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_6_io_in_psum = PE_Array_29_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_7_clock = clock;
  assign PE_Array_30_7_reset = reset;
  assign PE_Array_30_7_io_in_activate = PE_Array_30_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_7_io_in_weight = PE_Array_29_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_7_io_in_psum = PE_Array_29_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_8_clock = clock;
  assign PE_Array_30_8_reset = reset;
  assign PE_Array_30_8_io_in_activate = PE_Array_30_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_8_io_in_weight = PE_Array_29_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_8_io_in_psum = PE_Array_29_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_9_clock = clock;
  assign PE_Array_30_9_reset = reset;
  assign PE_Array_30_9_io_in_activate = PE_Array_30_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_9_io_in_weight = PE_Array_29_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_9_io_in_psum = PE_Array_29_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_10_clock = clock;
  assign PE_Array_30_10_reset = reset;
  assign PE_Array_30_10_io_in_activate = PE_Array_30_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_10_io_in_weight = PE_Array_29_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_10_io_in_psum = PE_Array_29_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_11_clock = clock;
  assign PE_Array_30_11_reset = reset;
  assign PE_Array_30_11_io_in_activate = PE_Array_30_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_11_io_in_weight = PE_Array_29_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_11_io_in_psum = PE_Array_29_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_12_clock = clock;
  assign PE_Array_30_12_reset = reset;
  assign PE_Array_30_12_io_in_activate = PE_Array_30_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_12_io_in_weight = PE_Array_29_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_12_io_in_psum = PE_Array_29_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_13_clock = clock;
  assign PE_Array_30_13_reset = reset;
  assign PE_Array_30_13_io_in_activate = PE_Array_30_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_13_io_in_weight = PE_Array_29_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_13_io_in_psum = PE_Array_29_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_14_clock = clock;
  assign PE_Array_30_14_reset = reset;
  assign PE_Array_30_14_io_in_activate = PE_Array_30_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_14_io_in_weight = PE_Array_29_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_14_io_in_psum = PE_Array_29_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_15_clock = clock;
  assign PE_Array_30_15_reset = reset;
  assign PE_Array_30_15_io_in_activate = PE_Array_30_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_15_io_in_weight = PE_Array_29_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_15_io_in_psum = PE_Array_29_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_16_clock = clock;
  assign PE_Array_30_16_reset = reset;
  assign PE_Array_30_16_io_in_activate = PE_Array_30_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_16_io_in_weight = PE_Array_29_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_16_io_in_psum = PE_Array_29_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_17_clock = clock;
  assign PE_Array_30_17_reset = reset;
  assign PE_Array_30_17_io_in_activate = PE_Array_30_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_17_io_in_weight = PE_Array_29_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_17_io_in_psum = PE_Array_29_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_18_clock = clock;
  assign PE_Array_30_18_reset = reset;
  assign PE_Array_30_18_io_in_activate = PE_Array_30_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_18_io_in_weight = PE_Array_29_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_18_io_in_psum = PE_Array_29_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_19_clock = clock;
  assign PE_Array_30_19_reset = reset;
  assign PE_Array_30_19_io_in_activate = PE_Array_30_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_19_io_in_weight = PE_Array_29_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_19_io_in_psum = PE_Array_29_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_20_clock = clock;
  assign PE_Array_30_20_reset = reset;
  assign PE_Array_30_20_io_in_activate = PE_Array_30_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_20_io_in_weight = PE_Array_29_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_20_io_in_psum = PE_Array_29_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_21_clock = clock;
  assign PE_Array_30_21_reset = reset;
  assign PE_Array_30_21_io_in_activate = PE_Array_30_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_21_io_in_weight = PE_Array_29_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_21_io_in_psum = PE_Array_29_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_22_clock = clock;
  assign PE_Array_30_22_reset = reset;
  assign PE_Array_30_22_io_in_activate = PE_Array_30_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_22_io_in_weight = PE_Array_29_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_22_io_in_psum = PE_Array_29_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_23_clock = clock;
  assign PE_Array_30_23_reset = reset;
  assign PE_Array_30_23_io_in_activate = PE_Array_30_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_23_io_in_weight = PE_Array_29_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_23_io_in_psum = PE_Array_29_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_24_clock = clock;
  assign PE_Array_30_24_reset = reset;
  assign PE_Array_30_24_io_in_activate = PE_Array_30_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_24_io_in_weight = PE_Array_29_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_24_io_in_psum = PE_Array_29_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_25_clock = clock;
  assign PE_Array_30_25_reset = reset;
  assign PE_Array_30_25_io_in_activate = PE_Array_30_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_25_io_in_weight = PE_Array_29_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_25_io_in_psum = PE_Array_29_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_26_clock = clock;
  assign PE_Array_30_26_reset = reset;
  assign PE_Array_30_26_io_in_activate = PE_Array_30_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_26_io_in_weight = PE_Array_29_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_26_io_in_psum = PE_Array_29_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_27_clock = clock;
  assign PE_Array_30_27_reset = reset;
  assign PE_Array_30_27_io_in_activate = PE_Array_30_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_27_io_in_weight = PE_Array_29_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_27_io_in_psum = PE_Array_29_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_28_clock = clock;
  assign PE_Array_30_28_reset = reset;
  assign PE_Array_30_28_io_in_activate = PE_Array_30_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_28_io_in_weight = PE_Array_29_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_28_io_in_psum = PE_Array_29_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_29_clock = clock;
  assign PE_Array_30_29_reset = reset;
  assign PE_Array_30_29_io_in_activate = PE_Array_30_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_29_io_in_weight = PE_Array_29_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_29_io_in_psum = PE_Array_29_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_30_clock = clock;
  assign PE_Array_30_30_reset = reset;
  assign PE_Array_30_30_io_in_activate = PE_Array_30_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_30_io_in_weight = PE_Array_29_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_30_io_in_psum = PE_Array_29_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_30_31_clock = clock;
  assign PE_Array_30_31_reset = reset;
  assign PE_Array_30_31_io_in_activate = PE_Array_30_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_30_31_io_in_weight = PE_Array_29_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_30_31_io_in_psum = PE_Array_29_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_30_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_30_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_0_clock = clock;
  assign PE_Array_31_0_reset = reset;
  assign PE_Array_31_0_io_in_activate = io_activate_31; // @[DataPath.scala 11:26]
  assign PE_Array_31_0_io_in_weight = PE_Array_30_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_0_io_in_psum = PE_Array_30_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_1_clock = clock;
  assign PE_Array_31_1_reset = reset;
  assign PE_Array_31_1_io_in_activate = PE_Array_31_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_1_io_in_weight = PE_Array_30_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_1_io_in_psum = PE_Array_30_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_2_clock = clock;
  assign PE_Array_31_2_reset = reset;
  assign PE_Array_31_2_io_in_activate = PE_Array_31_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_2_io_in_weight = PE_Array_30_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_2_io_in_psum = PE_Array_30_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_3_clock = clock;
  assign PE_Array_31_3_reset = reset;
  assign PE_Array_31_3_io_in_activate = PE_Array_31_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_3_io_in_weight = PE_Array_30_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_3_io_in_psum = PE_Array_30_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_4_clock = clock;
  assign PE_Array_31_4_reset = reset;
  assign PE_Array_31_4_io_in_activate = PE_Array_31_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_4_io_in_weight = PE_Array_30_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_4_io_in_psum = PE_Array_30_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_5_clock = clock;
  assign PE_Array_31_5_reset = reset;
  assign PE_Array_31_5_io_in_activate = PE_Array_31_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_5_io_in_weight = PE_Array_30_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_5_io_in_psum = PE_Array_30_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_6_clock = clock;
  assign PE_Array_31_6_reset = reset;
  assign PE_Array_31_6_io_in_activate = PE_Array_31_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_6_io_in_weight = PE_Array_30_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_6_io_in_psum = PE_Array_30_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_7_clock = clock;
  assign PE_Array_31_7_reset = reset;
  assign PE_Array_31_7_io_in_activate = PE_Array_31_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_7_io_in_weight = PE_Array_30_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_7_io_in_psum = PE_Array_30_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_8_clock = clock;
  assign PE_Array_31_8_reset = reset;
  assign PE_Array_31_8_io_in_activate = PE_Array_31_7_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_8_io_in_weight = PE_Array_30_8_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_8_io_in_psum = PE_Array_30_8_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_8_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_8_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_9_clock = clock;
  assign PE_Array_31_9_reset = reset;
  assign PE_Array_31_9_io_in_activate = PE_Array_31_8_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_9_io_in_weight = PE_Array_30_9_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_9_io_in_psum = PE_Array_30_9_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_9_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_9_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_10_clock = clock;
  assign PE_Array_31_10_reset = reset;
  assign PE_Array_31_10_io_in_activate = PE_Array_31_9_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_10_io_in_weight = PE_Array_30_10_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_10_io_in_psum = PE_Array_30_10_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_10_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_10_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_11_clock = clock;
  assign PE_Array_31_11_reset = reset;
  assign PE_Array_31_11_io_in_activate = PE_Array_31_10_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_11_io_in_weight = PE_Array_30_11_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_11_io_in_psum = PE_Array_30_11_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_11_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_11_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_12_clock = clock;
  assign PE_Array_31_12_reset = reset;
  assign PE_Array_31_12_io_in_activate = PE_Array_31_11_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_12_io_in_weight = PE_Array_30_12_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_12_io_in_psum = PE_Array_30_12_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_12_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_12_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_13_clock = clock;
  assign PE_Array_31_13_reset = reset;
  assign PE_Array_31_13_io_in_activate = PE_Array_31_12_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_13_io_in_weight = PE_Array_30_13_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_13_io_in_psum = PE_Array_30_13_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_13_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_13_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_14_clock = clock;
  assign PE_Array_31_14_reset = reset;
  assign PE_Array_31_14_io_in_activate = PE_Array_31_13_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_14_io_in_weight = PE_Array_30_14_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_14_io_in_psum = PE_Array_30_14_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_14_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_14_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_15_clock = clock;
  assign PE_Array_31_15_reset = reset;
  assign PE_Array_31_15_io_in_activate = PE_Array_31_14_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_15_io_in_weight = PE_Array_30_15_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_15_io_in_psum = PE_Array_30_15_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_15_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_15_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_16_clock = clock;
  assign PE_Array_31_16_reset = reset;
  assign PE_Array_31_16_io_in_activate = PE_Array_31_15_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_16_io_in_weight = PE_Array_30_16_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_16_io_in_psum = PE_Array_30_16_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_16_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_16_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_17_clock = clock;
  assign PE_Array_31_17_reset = reset;
  assign PE_Array_31_17_io_in_activate = PE_Array_31_16_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_17_io_in_weight = PE_Array_30_17_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_17_io_in_psum = PE_Array_30_17_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_17_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_17_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_18_clock = clock;
  assign PE_Array_31_18_reset = reset;
  assign PE_Array_31_18_io_in_activate = PE_Array_31_17_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_18_io_in_weight = PE_Array_30_18_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_18_io_in_psum = PE_Array_30_18_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_18_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_18_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_19_clock = clock;
  assign PE_Array_31_19_reset = reset;
  assign PE_Array_31_19_io_in_activate = PE_Array_31_18_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_19_io_in_weight = PE_Array_30_19_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_19_io_in_psum = PE_Array_30_19_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_19_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_19_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_20_clock = clock;
  assign PE_Array_31_20_reset = reset;
  assign PE_Array_31_20_io_in_activate = PE_Array_31_19_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_20_io_in_weight = PE_Array_30_20_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_20_io_in_psum = PE_Array_30_20_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_20_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_20_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_21_clock = clock;
  assign PE_Array_31_21_reset = reset;
  assign PE_Array_31_21_io_in_activate = PE_Array_31_20_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_21_io_in_weight = PE_Array_30_21_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_21_io_in_psum = PE_Array_30_21_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_21_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_21_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_22_clock = clock;
  assign PE_Array_31_22_reset = reset;
  assign PE_Array_31_22_io_in_activate = PE_Array_31_21_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_22_io_in_weight = PE_Array_30_22_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_22_io_in_psum = PE_Array_30_22_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_22_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_22_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_23_clock = clock;
  assign PE_Array_31_23_reset = reset;
  assign PE_Array_31_23_io_in_activate = PE_Array_31_22_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_23_io_in_weight = PE_Array_30_23_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_23_io_in_psum = PE_Array_30_23_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_23_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_23_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_24_clock = clock;
  assign PE_Array_31_24_reset = reset;
  assign PE_Array_31_24_io_in_activate = PE_Array_31_23_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_24_io_in_weight = PE_Array_30_24_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_24_io_in_psum = PE_Array_30_24_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_24_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_24_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_25_clock = clock;
  assign PE_Array_31_25_reset = reset;
  assign PE_Array_31_25_io_in_activate = PE_Array_31_24_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_25_io_in_weight = PE_Array_30_25_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_25_io_in_psum = PE_Array_30_25_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_25_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_25_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_26_clock = clock;
  assign PE_Array_31_26_reset = reset;
  assign PE_Array_31_26_io_in_activate = PE_Array_31_25_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_26_io_in_weight = PE_Array_30_26_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_26_io_in_psum = PE_Array_30_26_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_26_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_26_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_27_clock = clock;
  assign PE_Array_31_27_reset = reset;
  assign PE_Array_31_27_io_in_activate = PE_Array_31_26_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_27_io_in_weight = PE_Array_30_27_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_27_io_in_psum = PE_Array_30_27_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_27_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_27_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_28_clock = clock;
  assign PE_Array_31_28_reset = reset;
  assign PE_Array_31_28_io_in_activate = PE_Array_31_27_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_28_io_in_weight = PE_Array_30_28_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_28_io_in_psum = PE_Array_30_28_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_28_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_28_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_29_clock = clock;
  assign PE_Array_31_29_reset = reset;
  assign PE_Array_31_29_io_in_activate = PE_Array_31_28_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_29_io_in_weight = PE_Array_30_29_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_29_io_in_psum = PE_Array_30_29_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_29_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_29_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_30_clock = clock;
  assign PE_Array_31_30_reset = reset;
  assign PE_Array_31_30_io_in_activate = PE_Array_31_29_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_30_io_in_weight = PE_Array_30_30_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_30_io_in_psum = PE_Array_30_30_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_30_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_30_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_31_31_clock = clock;
  assign PE_Array_31_31_reset = reset;
  assign PE_Array_31_31_io_in_activate = PE_Array_31_30_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_31_31_io_in_weight = PE_Array_30_31_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_31_31_io_in_psum = PE_Array_30_31_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_31_31_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_31_31_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  always @(posedge clock) begin
    if (reset) begin // @[Systolic_Array.scala 52:29]
      flow_counter <= 7'h0; // @[Systolic_Array.scala 52:29]
    end else if (io_flow & flow_counter < 7'h5e) begin // @[Systolic_Array.scala 56:58]
      flow_counter <= _flow_counter_T_1; // @[Systolic_Array.scala 57:18]
    end else if (flow_counter == 7'h5e) begin // @[Systolic_Array.scala 58:53]
      flow_counter <= 7'h0; // @[Systolic_Array.scala 59:18]
    end
    if (reset) begin // @[Systolic_Array.scala 53:26]
      valid_reg <= 32'h0; // @[Systolic_Array.scala 53:26]
    end else if (io_flow & 7'h1f <= flow_counter & flow_counter < 7'h3f) begin // @[Systolic_Array.scala 65:96]
      valid_reg <= _valid_reg_T_1; // @[Systolic_Array.scala 66:15]
    end else if (io_flow & flow_counter >= 7'h3f) begin // @[Systolic_Array.scala 67:65]
      valid_reg <= _valid_reg_T_3; // @[Systolic_Array.scala 68:15]
    end else begin
      valid_reg <= 32'h0; // @[Systolic_Array.scala 70:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flow_counter = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
