module Activation_Buffer(
  input        clock,
  input        reset,
  input        io_wen,
  input        io_ren,
  input  [7:0] io_in_data_x_0,
  input  [7:0] io_in_data_x_1,
  input  [7:0] io_in_data_x_2,
  input  [7:0] io_in_data_x_3,
  input  [7:0] io_in_data_x_4,
  input  [7:0] io_in_data_x_5,
  input  [7:0] io_in_data_x_6,
  input  [7:0] io_in_data_x_7,
  input  [7:0] io_in_data_x_8,
  input  [7:0] io_in_data_x_9,
  input  [7:0] io_in_data_x_10,
  input  [7:0] io_in_data_x_11,
  input  [7:0] io_in_data_x_12,
  input  [7:0] io_in_data_x_13,
  input  [7:0] io_in_data_x_14,
  input  [7:0] io_in_data_x_15,
  input  [7:0] io_in_data_x_16,
  input  [7:0] io_in_data_x_17,
  input  [7:0] io_in_data_x_18,
  input  [7:0] io_in_data_x_19,
  input  [7:0] io_in_data_x_20,
  input  [7:0] io_in_data_x_21,
  input  [7:0] io_in_data_x_22,
  input  [7:0] io_in_data_x_23,
  input  [7:0] io_in_data_x_24,
  input  [7:0] io_in_data_x_25,
  input  [7:0] io_in_data_x_26,
  input  [7:0] io_in_data_x_27,
  input  [7:0] io_in_data_x_28,
  input  [7:0] io_in_data_x_29,
  input  [7:0] io_in_data_x_30,
  input  [7:0] io_in_data_x_31,
  input  [7:0] io_in_data_x_32,
  input  [7:0] io_in_data_x_33,
  input  [7:0] io_in_data_x_34,
  input  [7:0] io_in_data_x_35,
  input  [7:0] io_in_data_x_36,
  input  [7:0] io_in_data_x_37,
  input  [7:0] io_in_data_x_38,
  input  [7:0] io_in_data_x_39,
  input  [7:0] io_in_data_x_40,
  input  [7:0] io_in_data_x_41,
  input  [7:0] io_in_data_x_42,
  input  [7:0] io_in_data_x_43,
  input  [7:0] io_in_data_x_44,
  input  [7:0] io_in_data_x_45,
  input  [7:0] io_in_data_x_46,
  input  [7:0] io_in_data_x_47,
  input  [7:0] io_in_data_x_48,
  input  [7:0] io_in_data_x_49,
  input  [7:0] io_in_data_x_50,
  input  [7:0] io_in_data_x_51,
  input  [7:0] io_in_data_x_52,
  input  [7:0] io_in_data_x_53,
  input  [7:0] io_in_data_x_54,
  input  [7:0] io_in_data_x_55,
  input  [7:0] io_in_data_x_56,
  input  [7:0] io_in_data_x_57,
  input  [7:0] io_in_data_x_58,
  input  [7:0] io_in_data_x_59,
  input  [7:0] io_in_data_x_60,
  input  [7:0] io_in_data_x_61,
  input  [7:0] io_in_data_x_62,
  input  [7:0] io_in_data_x_63,
  output [7:0] io_out_activate_0,
  output [7:0] io_out_activate_1,
  output [7:0] io_out_activate_2,
  output [7:0] io_out_activate_3,
  output [7:0] io_out_activate_4,
  output [7:0] io_out_activate_5,
  output [7:0] io_out_activate_6,
  output [7:0] io_out_activate_7,
  output       io_out_flow,
  output       io_isfull,
  output       io_isempty,
  output       io_isdone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] buffer_0_0; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_1; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_2; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_3; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_4; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_5; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_6; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_7; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_8; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_9; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_10; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_11; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_12; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_13; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_14; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_15; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_16; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_17; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_18; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_19; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_20; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_21; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_22; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_23; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_24; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_25; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_26; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_27; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_28; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_29; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_30; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_31; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_32; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_33; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_34; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_35; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_36; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_37; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_38; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_39; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_40; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_41; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_42; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_43; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_44; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_45; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_46; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_47; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_48; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_49; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_50; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_51; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_52; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_53; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_54; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_55; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_56; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_57; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_58; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_59; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_60; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_61; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_62; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_0_63; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_0; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_1; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_2; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_3; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_4; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_5; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_6; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_7; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_8; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_9; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_10; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_11; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_12; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_13; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_14; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_15; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_16; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_17; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_18; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_19; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_20; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_21; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_22; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_23; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_24; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_25; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_26; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_27; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_28; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_29; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_30; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_31; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_32; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_33; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_34; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_35; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_36; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_37; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_38; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_39; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_40; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_41; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_42; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_43; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_44; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_45; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_46; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_47; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_48; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_49; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_50; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_51; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_52; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_53; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_54; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_55; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_56; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_57; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_58; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_59; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_60; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_61; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_62; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_1_63; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_0; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_1; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_2; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_3; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_4; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_5; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_6; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_7; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_8; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_9; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_10; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_11; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_12; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_13; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_14; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_15; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_16; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_17; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_18; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_19; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_20; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_21; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_22; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_23; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_24; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_25; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_26; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_27; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_28; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_29; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_30; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_31; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_32; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_33; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_34; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_35; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_36; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_37; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_38; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_39; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_40; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_41; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_42; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_43; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_44; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_45; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_46; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_47; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_48; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_49; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_50; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_51; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_52; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_53; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_54; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_55; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_56; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_57; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_58; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_59; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_60; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_61; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_62; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_2_63; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_0; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_1; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_2; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_3; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_4; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_5; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_6; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_7; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_8; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_9; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_10; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_11; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_12; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_13; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_14; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_15; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_16; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_17; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_18; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_19; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_20; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_21; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_22; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_23; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_24; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_25; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_26; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_27; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_28; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_29; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_30; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_31; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_32; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_33; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_34; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_35; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_36; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_37; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_38; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_39; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_40; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_41; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_42; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_43; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_44; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_45; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_46; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_47; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_48; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_49; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_50; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_51; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_52; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_53; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_54; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_55; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_56; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_57; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_58; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_59; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_60; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_61; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_62; // @[Activation_Buffer.scala 24:23]
  reg [7:0] buffer_3_63; // @[Activation_Buffer.scala 24:23]
  reg [2:0] read_ptr; // @[Activation_Buffer.scala 27:25]
  reg [2:0] write_ptr; // @[Activation_Buffer.scala 28:26]
  wire  _full_T_2 = read_ptr[1:0] == write_ptr[1:0]; // @[Activation_Buffer.scala 33:44]
  wire  full = read_ptr[1:0] == write_ptr[1:0] & read_ptr[2] != write_ptr[2]; // @[Activation_Buffer.scala 33:82]
  wire  empty = _full_T_2 & read_ptr[2] == write_ptr[2]; // @[Activation_Buffer.scala 34:83]
  wire  _T_1 = io_wen & ~full; // @[Activation_Buffer.scala 39:15]
  wire [2:0] _write_ptr_T_1 = write_ptr + 3'h1; // @[Activation_Buffer.scala 40:28]
  reg [4:0] flow_ptr; // @[Activation_Buffer.scala 55:25]
  wire [4:0] _flow_ptr_T_1 = flow_ptr + 5'h1; // @[Activation_Buffer.scala 58:26]
  wire  _T_70 = flow_ptr == 5'h16; // @[Activation_Buffer.scala 59:23]
  wire  _T_71 = flow_ptr != 5'h0; // @[Activation_Buffer.scala 61:23]
  wire [5:0] _io_out_activate_0_T_1 = {{1'd0}, flow_ptr}; // @[Activation_Buffer.scala 76:88]
  wire [4:0] _io_out_activate_0_T_4 = _io_out_activate_0_T_1[4:0] - 5'h1; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_518 = 2'h0 == read_ptr[1:0] & 5'h1 == _io_out_activate_0_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_519 = 2'h0 == read_ptr[1:0] & 5'h2 == _io_out_activate_0_T_4 ? buffer_0_2 : _GEN_518; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_520 = 2'h0 == read_ptr[1:0] & 5'h3 == _io_out_activate_0_T_4 ? buffer_0_3 : _GEN_519; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_521 = 2'h0 == read_ptr[1:0] & 5'h4 == _io_out_activate_0_T_4 ? buffer_0_4 : _GEN_520; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_522 = 2'h0 == read_ptr[1:0] & 5'h5 == _io_out_activate_0_T_4 ? buffer_0_5 : _GEN_521; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_523 = 2'h0 == read_ptr[1:0] & 5'h6 == _io_out_activate_0_T_4 ? buffer_0_6 : _GEN_522; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_524 = 2'h0 == read_ptr[1:0] & 5'h7 == _io_out_activate_0_T_4 ? buffer_0_7 : _GEN_523; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_525 = 2'h0 == read_ptr[1:0] & 5'h8 == _io_out_activate_0_T_4 ? buffer_0_8 : _GEN_524; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_526 = 2'h0 == read_ptr[1:0] & 5'h9 == _io_out_activate_0_T_4 ? buffer_0_9 : _GEN_525; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_527 = 2'h0 == read_ptr[1:0] & 5'ha == _io_out_activate_0_T_4 ? buffer_0_10 : _GEN_526; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_528 = 2'h0 == read_ptr[1:0] & 5'hb == _io_out_activate_0_T_4 ? buffer_0_11 : _GEN_527; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_529 = 2'h0 == read_ptr[1:0] & 5'hc == _io_out_activate_0_T_4 ? buffer_0_12 : _GEN_528; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_530 = 2'h0 == read_ptr[1:0] & 5'hd == _io_out_activate_0_T_4 ? buffer_0_13 : _GEN_529; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_531 = 2'h0 == read_ptr[1:0] & 5'he == _io_out_activate_0_T_4 ? buffer_0_14 : _GEN_530; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_532 = 2'h0 == read_ptr[1:0] & 5'hf == _io_out_activate_0_T_4 ? buffer_0_15 : _GEN_531; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_533 = 2'h0 == read_ptr[1:0] & 5'h10 == _io_out_activate_0_T_4 ? buffer_0_16 : _GEN_532; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_534 = 2'h0 == read_ptr[1:0] & 5'h11 == _io_out_activate_0_T_4 ? buffer_0_17 : _GEN_533; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_535 = 2'h0 == read_ptr[1:0] & 5'h12 == _io_out_activate_0_T_4 ? buffer_0_18 : _GEN_534; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_536 = 2'h0 == read_ptr[1:0] & 5'h13 == _io_out_activate_0_T_4 ? buffer_0_19 : _GEN_535; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_537 = 2'h0 == read_ptr[1:0] & 5'h14 == _io_out_activate_0_T_4 ? buffer_0_20 : _GEN_536; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_538 = 2'h0 == read_ptr[1:0] & 5'h15 == _io_out_activate_0_T_4 ? buffer_0_21 : _GEN_537; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_539 = 2'h0 == read_ptr[1:0] & 5'h16 == _io_out_activate_0_T_4 ? buffer_0_22 : _GEN_538; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_540 = 2'h0 == read_ptr[1:0] & 5'h17 == _io_out_activate_0_T_4 ? buffer_0_23 : _GEN_539; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_541 = 2'h0 == read_ptr[1:0] & 5'h18 == _io_out_activate_0_T_4 ? buffer_0_24 : _GEN_540; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_542 = 2'h0 == read_ptr[1:0] & 5'h19 == _io_out_activate_0_T_4 ? buffer_0_25 : _GEN_541; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_543 = 2'h0 == read_ptr[1:0] & 5'h1a == _io_out_activate_0_T_4 ? buffer_0_26 : _GEN_542; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_544 = 2'h0 == read_ptr[1:0] & 5'h1b == _io_out_activate_0_T_4 ? buffer_0_27 : _GEN_543; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_545 = 2'h0 == read_ptr[1:0] & 5'h1c == _io_out_activate_0_T_4 ? buffer_0_28 : _GEN_544; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_546 = 2'h0 == read_ptr[1:0] & 5'h1d == _io_out_activate_0_T_4 ? buffer_0_29 : _GEN_545; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_547 = 2'h0 == read_ptr[1:0] & 5'h1e == _io_out_activate_0_T_4 ? buffer_0_30 : _GEN_546; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_548 = 2'h0 == read_ptr[1:0] & 5'h1f == _io_out_activate_0_T_4 ? buffer_0_31 : _GEN_547; // @[Activation_Buffer.scala 76:{28,28}]
  wire [5:0] _GEN_2645 = {{1'd0}, _io_out_activate_0_T_4}; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_549 = 2'h0 == read_ptr[1:0] & 6'h20 == _GEN_2645 ? buffer_0_32 : _GEN_548; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_550 = 2'h0 == read_ptr[1:0] & 6'h21 == _GEN_2645 ? buffer_0_33 : _GEN_549; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_551 = 2'h0 == read_ptr[1:0] & 6'h22 == _GEN_2645 ? buffer_0_34 : _GEN_550; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_552 = 2'h0 == read_ptr[1:0] & 6'h23 == _GEN_2645 ? buffer_0_35 : _GEN_551; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_553 = 2'h0 == read_ptr[1:0] & 6'h24 == _GEN_2645 ? buffer_0_36 : _GEN_552; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_554 = 2'h0 == read_ptr[1:0] & 6'h25 == _GEN_2645 ? buffer_0_37 : _GEN_553; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_555 = 2'h0 == read_ptr[1:0] & 6'h26 == _GEN_2645 ? buffer_0_38 : _GEN_554; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_556 = 2'h0 == read_ptr[1:0] & 6'h27 == _GEN_2645 ? buffer_0_39 : _GEN_555; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_557 = 2'h0 == read_ptr[1:0] & 6'h28 == _GEN_2645 ? buffer_0_40 : _GEN_556; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_558 = 2'h0 == read_ptr[1:0] & 6'h29 == _GEN_2645 ? buffer_0_41 : _GEN_557; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_559 = 2'h0 == read_ptr[1:0] & 6'h2a == _GEN_2645 ? buffer_0_42 : _GEN_558; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_560 = 2'h0 == read_ptr[1:0] & 6'h2b == _GEN_2645 ? buffer_0_43 : _GEN_559; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_561 = 2'h0 == read_ptr[1:0] & 6'h2c == _GEN_2645 ? buffer_0_44 : _GEN_560; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_562 = 2'h0 == read_ptr[1:0] & 6'h2d == _GEN_2645 ? buffer_0_45 : _GEN_561; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_563 = 2'h0 == read_ptr[1:0] & 6'h2e == _GEN_2645 ? buffer_0_46 : _GEN_562; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_564 = 2'h0 == read_ptr[1:0] & 6'h2f == _GEN_2645 ? buffer_0_47 : _GEN_563; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_565 = 2'h0 == read_ptr[1:0] & 6'h30 == _GEN_2645 ? buffer_0_48 : _GEN_564; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_566 = 2'h0 == read_ptr[1:0] & 6'h31 == _GEN_2645 ? buffer_0_49 : _GEN_565; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_567 = 2'h0 == read_ptr[1:0] & 6'h32 == _GEN_2645 ? buffer_0_50 : _GEN_566; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_568 = 2'h0 == read_ptr[1:0] & 6'h33 == _GEN_2645 ? buffer_0_51 : _GEN_567; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_569 = 2'h0 == read_ptr[1:0] & 6'h34 == _GEN_2645 ? buffer_0_52 : _GEN_568; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_570 = 2'h0 == read_ptr[1:0] & 6'h35 == _GEN_2645 ? buffer_0_53 : _GEN_569; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_571 = 2'h0 == read_ptr[1:0] & 6'h36 == _GEN_2645 ? buffer_0_54 : _GEN_570; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_572 = 2'h0 == read_ptr[1:0] & 6'h37 == _GEN_2645 ? buffer_0_55 : _GEN_571; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_573 = 2'h0 == read_ptr[1:0] & 6'h38 == _GEN_2645 ? buffer_0_56 : _GEN_572; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_574 = 2'h0 == read_ptr[1:0] & 6'h39 == _GEN_2645 ? buffer_0_57 : _GEN_573; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_575 = 2'h0 == read_ptr[1:0] & 6'h3a == _GEN_2645 ? buffer_0_58 : _GEN_574; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_576 = 2'h0 == read_ptr[1:0] & 6'h3b == _GEN_2645 ? buffer_0_59 : _GEN_575; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_577 = 2'h0 == read_ptr[1:0] & 6'h3c == _GEN_2645 ? buffer_0_60 : _GEN_576; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_578 = 2'h0 == read_ptr[1:0] & 6'h3d == _GEN_2645 ? buffer_0_61 : _GEN_577; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_579 = 2'h0 == read_ptr[1:0] & 6'h3e == _GEN_2645 ? buffer_0_62 : _GEN_578; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_580 = 2'h0 == read_ptr[1:0] & 6'h3f == _GEN_2645 ? buffer_0_63 : _GEN_579; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_581 = 2'h1 == read_ptr[1:0] & 5'h0 == _io_out_activate_0_T_4 ? buffer_1_0 : _GEN_580; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_582 = 2'h1 == read_ptr[1:0] & 5'h1 == _io_out_activate_0_T_4 ? buffer_1_1 : _GEN_581; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_583 = 2'h1 == read_ptr[1:0] & 5'h2 == _io_out_activate_0_T_4 ? buffer_1_2 : _GEN_582; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_584 = 2'h1 == read_ptr[1:0] & 5'h3 == _io_out_activate_0_T_4 ? buffer_1_3 : _GEN_583; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_585 = 2'h1 == read_ptr[1:0] & 5'h4 == _io_out_activate_0_T_4 ? buffer_1_4 : _GEN_584; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_586 = 2'h1 == read_ptr[1:0] & 5'h5 == _io_out_activate_0_T_4 ? buffer_1_5 : _GEN_585; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_587 = 2'h1 == read_ptr[1:0] & 5'h6 == _io_out_activate_0_T_4 ? buffer_1_6 : _GEN_586; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_588 = 2'h1 == read_ptr[1:0] & 5'h7 == _io_out_activate_0_T_4 ? buffer_1_7 : _GEN_587; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_589 = 2'h1 == read_ptr[1:0] & 5'h8 == _io_out_activate_0_T_4 ? buffer_1_8 : _GEN_588; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_590 = 2'h1 == read_ptr[1:0] & 5'h9 == _io_out_activate_0_T_4 ? buffer_1_9 : _GEN_589; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_591 = 2'h1 == read_ptr[1:0] & 5'ha == _io_out_activate_0_T_4 ? buffer_1_10 : _GEN_590; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_592 = 2'h1 == read_ptr[1:0] & 5'hb == _io_out_activate_0_T_4 ? buffer_1_11 : _GEN_591; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_593 = 2'h1 == read_ptr[1:0] & 5'hc == _io_out_activate_0_T_4 ? buffer_1_12 : _GEN_592; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_594 = 2'h1 == read_ptr[1:0] & 5'hd == _io_out_activate_0_T_4 ? buffer_1_13 : _GEN_593; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_595 = 2'h1 == read_ptr[1:0] & 5'he == _io_out_activate_0_T_4 ? buffer_1_14 : _GEN_594; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_596 = 2'h1 == read_ptr[1:0] & 5'hf == _io_out_activate_0_T_4 ? buffer_1_15 : _GEN_595; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_597 = 2'h1 == read_ptr[1:0] & 5'h10 == _io_out_activate_0_T_4 ? buffer_1_16 : _GEN_596; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_598 = 2'h1 == read_ptr[1:0] & 5'h11 == _io_out_activate_0_T_4 ? buffer_1_17 : _GEN_597; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_599 = 2'h1 == read_ptr[1:0] & 5'h12 == _io_out_activate_0_T_4 ? buffer_1_18 : _GEN_598; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_600 = 2'h1 == read_ptr[1:0] & 5'h13 == _io_out_activate_0_T_4 ? buffer_1_19 : _GEN_599; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_601 = 2'h1 == read_ptr[1:0] & 5'h14 == _io_out_activate_0_T_4 ? buffer_1_20 : _GEN_600; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_602 = 2'h1 == read_ptr[1:0] & 5'h15 == _io_out_activate_0_T_4 ? buffer_1_21 : _GEN_601; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_603 = 2'h1 == read_ptr[1:0] & 5'h16 == _io_out_activate_0_T_4 ? buffer_1_22 : _GEN_602; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_604 = 2'h1 == read_ptr[1:0] & 5'h17 == _io_out_activate_0_T_4 ? buffer_1_23 : _GEN_603; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_605 = 2'h1 == read_ptr[1:0] & 5'h18 == _io_out_activate_0_T_4 ? buffer_1_24 : _GEN_604; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_606 = 2'h1 == read_ptr[1:0] & 5'h19 == _io_out_activate_0_T_4 ? buffer_1_25 : _GEN_605; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_607 = 2'h1 == read_ptr[1:0] & 5'h1a == _io_out_activate_0_T_4 ? buffer_1_26 : _GEN_606; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_608 = 2'h1 == read_ptr[1:0] & 5'h1b == _io_out_activate_0_T_4 ? buffer_1_27 : _GEN_607; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_609 = 2'h1 == read_ptr[1:0] & 5'h1c == _io_out_activate_0_T_4 ? buffer_1_28 : _GEN_608; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_610 = 2'h1 == read_ptr[1:0] & 5'h1d == _io_out_activate_0_T_4 ? buffer_1_29 : _GEN_609; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_611 = 2'h1 == read_ptr[1:0] & 5'h1e == _io_out_activate_0_T_4 ? buffer_1_30 : _GEN_610; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_612 = 2'h1 == read_ptr[1:0] & 5'h1f == _io_out_activate_0_T_4 ? buffer_1_31 : _GEN_611; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_613 = 2'h1 == read_ptr[1:0] & 6'h20 == _GEN_2645 ? buffer_1_32 : _GEN_612; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_614 = 2'h1 == read_ptr[1:0] & 6'h21 == _GEN_2645 ? buffer_1_33 : _GEN_613; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_615 = 2'h1 == read_ptr[1:0] & 6'h22 == _GEN_2645 ? buffer_1_34 : _GEN_614; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_616 = 2'h1 == read_ptr[1:0] & 6'h23 == _GEN_2645 ? buffer_1_35 : _GEN_615; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_617 = 2'h1 == read_ptr[1:0] & 6'h24 == _GEN_2645 ? buffer_1_36 : _GEN_616; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_618 = 2'h1 == read_ptr[1:0] & 6'h25 == _GEN_2645 ? buffer_1_37 : _GEN_617; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_619 = 2'h1 == read_ptr[1:0] & 6'h26 == _GEN_2645 ? buffer_1_38 : _GEN_618; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_620 = 2'h1 == read_ptr[1:0] & 6'h27 == _GEN_2645 ? buffer_1_39 : _GEN_619; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_621 = 2'h1 == read_ptr[1:0] & 6'h28 == _GEN_2645 ? buffer_1_40 : _GEN_620; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_622 = 2'h1 == read_ptr[1:0] & 6'h29 == _GEN_2645 ? buffer_1_41 : _GEN_621; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_623 = 2'h1 == read_ptr[1:0] & 6'h2a == _GEN_2645 ? buffer_1_42 : _GEN_622; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_624 = 2'h1 == read_ptr[1:0] & 6'h2b == _GEN_2645 ? buffer_1_43 : _GEN_623; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_625 = 2'h1 == read_ptr[1:0] & 6'h2c == _GEN_2645 ? buffer_1_44 : _GEN_624; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_626 = 2'h1 == read_ptr[1:0] & 6'h2d == _GEN_2645 ? buffer_1_45 : _GEN_625; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_627 = 2'h1 == read_ptr[1:0] & 6'h2e == _GEN_2645 ? buffer_1_46 : _GEN_626; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_628 = 2'h1 == read_ptr[1:0] & 6'h2f == _GEN_2645 ? buffer_1_47 : _GEN_627; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_629 = 2'h1 == read_ptr[1:0] & 6'h30 == _GEN_2645 ? buffer_1_48 : _GEN_628; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_630 = 2'h1 == read_ptr[1:0] & 6'h31 == _GEN_2645 ? buffer_1_49 : _GEN_629; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_631 = 2'h1 == read_ptr[1:0] & 6'h32 == _GEN_2645 ? buffer_1_50 : _GEN_630; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_632 = 2'h1 == read_ptr[1:0] & 6'h33 == _GEN_2645 ? buffer_1_51 : _GEN_631; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_633 = 2'h1 == read_ptr[1:0] & 6'h34 == _GEN_2645 ? buffer_1_52 : _GEN_632; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_634 = 2'h1 == read_ptr[1:0] & 6'h35 == _GEN_2645 ? buffer_1_53 : _GEN_633; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_635 = 2'h1 == read_ptr[1:0] & 6'h36 == _GEN_2645 ? buffer_1_54 : _GEN_634; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_636 = 2'h1 == read_ptr[1:0] & 6'h37 == _GEN_2645 ? buffer_1_55 : _GEN_635; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_637 = 2'h1 == read_ptr[1:0] & 6'h38 == _GEN_2645 ? buffer_1_56 : _GEN_636; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_638 = 2'h1 == read_ptr[1:0] & 6'h39 == _GEN_2645 ? buffer_1_57 : _GEN_637; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_639 = 2'h1 == read_ptr[1:0] & 6'h3a == _GEN_2645 ? buffer_1_58 : _GEN_638; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_640 = 2'h1 == read_ptr[1:0] & 6'h3b == _GEN_2645 ? buffer_1_59 : _GEN_639; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_641 = 2'h1 == read_ptr[1:0] & 6'h3c == _GEN_2645 ? buffer_1_60 : _GEN_640; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_642 = 2'h1 == read_ptr[1:0] & 6'h3d == _GEN_2645 ? buffer_1_61 : _GEN_641; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_643 = 2'h1 == read_ptr[1:0] & 6'h3e == _GEN_2645 ? buffer_1_62 : _GEN_642; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_644 = 2'h1 == read_ptr[1:0] & 6'h3f == _GEN_2645 ? buffer_1_63 : _GEN_643; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_645 = 2'h2 == read_ptr[1:0] & 5'h0 == _io_out_activate_0_T_4 ? buffer_2_0 : _GEN_644; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_646 = 2'h2 == read_ptr[1:0] & 5'h1 == _io_out_activate_0_T_4 ? buffer_2_1 : _GEN_645; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_647 = 2'h2 == read_ptr[1:0] & 5'h2 == _io_out_activate_0_T_4 ? buffer_2_2 : _GEN_646; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_648 = 2'h2 == read_ptr[1:0] & 5'h3 == _io_out_activate_0_T_4 ? buffer_2_3 : _GEN_647; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_649 = 2'h2 == read_ptr[1:0] & 5'h4 == _io_out_activate_0_T_4 ? buffer_2_4 : _GEN_648; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_650 = 2'h2 == read_ptr[1:0] & 5'h5 == _io_out_activate_0_T_4 ? buffer_2_5 : _GEN_649; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_651 = 2'h2 == read_ptr[1:0] & 5'h6 == _io_out_activate_0_T_4 ? buffer_2_6 : _GEN_650; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_652 = 2'h2 == read_ptr[1:0] & 5'h7 == _io_out_activate_0_T_4 ? buffer_2_7 : _GEN_651; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_653 = 2'h2 == read_ptr[1:0] & 5'h8 == _io_out_activate_0_T_4 ? buffer_2_8 : _GEN_652; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_654 = 2'h2 == read_ptr[1:0] & 5'h9 == _io_out_activate_0_T_4 ? buffer_2_9 : _GEN_653; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_655 = 2'h2 == read_ptr[1:0] & 5'ha == _io_out_activate_0_T_4 ? buffer_2_10 : _GEN_654; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_656 = 2'h2 == read_ptr[1:0] & 5'hb == _io_out_activate_0_T_4 ? buffer_2_11 : _GEN_655; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_657 = 2'h2 == read_ptr[1:0] & 5'hc == _io_out_activate_0_T_4 ? buffer_2_12 : _GEN_656; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_658 = 2'h2 == read_ptr[1:0] & 5'hd == _io_out_activate_0_T_4 ? buffer_2_13 : _GEN_657; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_659 = 2'h2 == read_ptr[1:0] & 5'he == _io_out_activate_0_T_4 ? buffer_2_14 : _GEN_658; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_660 = 2'h2 == read_ptr[1:0] & 5'hf == _io_out_activate_0_T_4 ? buffer_2_15 : _GEN_659; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_661 = 2'h2 == read_ptr[1:0] & 5'h10 == _io_out_activate_0_T_4 ? buffer_2_16 : _GEN_660; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_662 = 2'h2 == read_ptr[1:0] & 5'h11 == _io_out_activate_0_T_4 ? buffer_2_17 : _GEN_661; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_663 = 2'h2 == read_ptr[1:0] & 5'h12 == _io_out_activate_0_T_4 ? buffer_2_18 : _GEN_662; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_664 = 2'h2 == read_ptr[1:0] & 5'h13 == _io_out_activate_0_T_4 ? buffer_2_19 : _GEN_663; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_665 = 2'h2 == read_ptr[1:0] & 5'h14 == _io_out_activate_0_T_4 ? buffer_2_20 : _GEN_664; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_666 = 2'h2 == read_ptr[1:0] & 5'h15 == _io_out_activate_0_T_4 ? buffer_2_21 : _GEN_665; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_667 = 2'h2 == read_ptr[1:0] & 5'h16 == _io_out_activate_0_T_4 ? buffer_2_22 : _GEN_666; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_668 = 2'h2 == read_ptr[1:0] & 5'h17 == _io_out_activate_0_T_4 ? buffer_2_23 : _GEN_667; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_669 = 2'h2 == read_ptr[1:0] & 5'h18 == _io_out_activate_0_T_4 ? buffer_2_24 : _GEN_668; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_670 = 2'h2 == read_ptr[1:0] & 5'h19 == _io_out_activate_0_T_4 ? buffer_2_25 : _GEN_669; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_671 = 2'h2 == read_ptr[1:0] & 5'h1a == _io_out_activate_0_T_4 ? buffer_2_26 : _GEN_670; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_672 = 2'h2 == read_ptr[1:0] & 5'h1b == _io_out_activate_0_T_4 ? buffer_2_27 : _GEN_671; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_673 = 2'h2 == read_ptr[1:0] & 5'h1c == _io_out_activate_0_T_4 ? buffer_2_28 : _GEN_672; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_674 = 2'h2 == read_ptr[1:0] & 5'h1d == _io_out_activate_0_T_4 ? buffer_2_29 : _GEN_673; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_675 = 2'h2 == read_ptr[1:0] & 5'h1e == _io_out_activate_0_T_4 ? buffer_2_30 : _GEN_674; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_676 = 2'h2 == read_ptr[1:0] & 5'h1f == _io_out_activate_0_T_4 ? buffer_2_31 : _GEN_675; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_677 = 2'h2 == read_ptr[1:0] & 6'h20 == _GEN_2645 ? buffer_2_32 : _GEN_676; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_678 = 2'h2 == read_ptr[1:0] & 6'h21 == _GEN_2645 ? buffer_2_33 : _GEN_677; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_679 = 2'h2 == read_ptr[1:0] & 6'h22 == _GEN_2645 ? buffer_2_34 : _GEN_678; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_680 = 2'h2 == read_ptr[1:0] & 6'h23 == _GEN_2645 ? buffer_2_35 : _GEN_679; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_681 = 2'h2 == read_ptr[1:0] & 6'h24 == _GEN_2645 ? buffer_2_36 : _GEN_680; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_682 = 2'h2 == read_ptr[1:0] & 6'h25 == _GEN_2645 ? buffer_2_37 : _GEN_681; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_683 = 2'h2 == read_ptr[1:0] & 6'h26 == _GEN_2645 ? buffer_2_38 : _GEN_682; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_684 = 2'h2 == read_ptr[1:0] & 6'h27 == _GEN_2645 ? buffer_2_39 : _GEN_683; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_685 = 2'h2 == read_ptr[1:0] & 6'h28 == _GEN_2645 ? buffer_2_40 : _GEN_684; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_686 = 2'h2 == read_ptr[1:0] & 6'h29 == _GEN_2645 ? buffer_2_41 : _GEN_685; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_687 = 2'h2 == read_ptr[1:0] & 6'h2a == _GEN_2645 ? buffer_2_42 : _GEN_686; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_688 = 2'h2 == read_ptr[1:0] & 6'h2b == _GEN_2645 ? buffer_2_43 : _GEN_687; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_689 = 2'h2 == read_ptr[1:0] & 6'h2c == _GEN_2645 ? buffer_2_44 : _GEN_688; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_690 = 2'h2 == read_ptr[1:0] & 6'h2d == _GEN_2645 ? buffer_2_45 : _GEN_689; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_691 = 2'h2 == read_ptr[1:0] & 6'h2e == _GEN_2645 ? buffer_2_46 : _GEN_690; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_692 = 2'h2 == read_ptr[1:0] & 6'h2f == _GEN_2645 ? buffer_2_47 : _GEN_691; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_693 = 2'h2 == read_ptr[1:0] & 6'h30 == _GEN_2645 ? buffer_2_48 : _GEN_692; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_694 = 2'h2 == read_ptr[1:0] & 6'h31 == _GEN_2645 ? buffer_2_49 : _GEN_693; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_695 = 2'h2 == read_ptr[1:0] & 6'h32 == _GEN_2645 ? buffer_2_50 : _GEN_694; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_696 = 2'h2 == read_ptr[1:0] & 6'h33 == _GEN_2645 ? buffer_2_51 : _GEN_695; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_697 = 2'h2 == read_ptr[1:0] & 6'h34 == _GEN_2645 ? buffer_2_52 : _GEN_696; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_698 = 2'h2 == read_ptr[1:0] & 6'h35 == _GEN_2645 ? buffer_2_53 : _GEN_697; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_699 = 2'h2 == read_ptr[1:0] & 6'h36 == _GEN_2645 ? buffer_2_54 : _GEN_698; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_700 = 2'h2 == read_ptr[1:0] & 6'h37 == _GEN_2645 ? buffer_2_55 : _GEN_699; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_701 = 2'h2 == read_ptr[1:0] & 6'h38 == _GEN_2645 ? buffer_2_56 : _GEN_700; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_702 = 2'h2 == read_ptr[1:0] & 6'h39 == _GEN_2645 ? buffer_2_57 : _GEN_701; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_703 = 2'h2 == read_ptr[1:0] & 6'h3a == _GEN_2645 ? buffer_2_58 : _GEN_702; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_704 = 2'h2 == read_ptr[1:0] & 6'h3b == _GEN_2645 ? buffer_2_59 : _GEN_703; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_705 = 2'h2 == read_ptr[1:0] & 6'h3c == _GEN_2645 ? buffer_2_60 : _GEN_704; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_706 = 2'h2 == read_ptr[1:0] & 6'h3d == _GEN_2645 ? buffer_2_61 : _GEN_705; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_707 = 2'h2 == read_ptr[1:0] & 6'h3e == _GEN_2645 ? buffer_2_62 : _GEN_706; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_708 = 2'h2 == read_ptr[1:0] & 6'h3f == _GEN_2645 ? buffer_2_63 : _GEN_707; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_709 = 2'h3 == read_ptr[1:0] & 5'h0 == _io_out_activate_0_T_4 ? buffer_3_0 : _GEN_708; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_710 = 2'h3 == read_ptr[1:0] & 5'h1 == _io_out_activate_0_T_4 ? buffer_3_1 : _GEN_709; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_711 = 2'h3 == read_ptr[1:0] & 5'h2 == _io_out_activate_0_T_4 ? buffer_3_2 : _GEN_710; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_712 = 2'h3 == read_ptr[1:0] & 5'h3 == _io_out_activate_0_T_4 ? buffer_3_3 : _GEN_711; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_713 = 2'h3 == read_ptr[1:0] & 5'h4 == _io_out_activate_0_T_4 ? buffer_3_4 : _GEN_712; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_714 = 2'h3 == read_ptr[1:0] & 5'h5 == _io_out_activate_0_T_4 ? buffer_3_5 : _GEN_713; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_715 = 2'h3 == read_ptr[1:0] & 5'h6 == _io_out_activate_0_T_4 ? buffer_3_6 : _GEN_714; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_716 = 2'h3 == read_ptr[1:0] & 5'h7 == _io_out_activate_0_T_4 ? buffer_3_7 : _GEN_715; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_717 = 2'h3 == read_ptr[1:0] & 5'h8 == _io_out_activate_0_T_4 ? buffer_3_8 : _GEN_716; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_718 = 2'h3 == read_ptr[1:0] & 5'h9 == _io_out_activate_0_T_4 ? buffer_3_9 : _GEN_717; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_719 = 2'h3 == read_ptr[1:0] & 5'ha == _io_out_activate_0_T_4 ? buffer_3_10 : _GEN_718; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_720 = 2'h3 == read_ptr[1:0] & 5'hb == _io_out_activate_0_T_4 ? buffer_3_11 : _GEN_719; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_721 = 2'h3 == read_ptr[1:0] & 5'hc == _io_out_activate_0_T_4 ? buffer_3_12 : _GEN_720; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_722 = 2'h3 == read_ptr[1:0] & 5'hd == _io_out_activate_0_T_4 ? buffer_3_13 : _GEN_721; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_723 = 2'h3 == read_ptr[1:0] & 5'he == _io_out_activate_0_T_4 ? buffer_3_14 : _GEN_722; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_724 = 2'h3 == read_ptr[1:0] & 5'hf == _io_out_activate_0_T_4 ? buffer_3_15 : _GEN_723; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_725 = 2'h3 == read_ptr[1:0] & 5'h10 == _io_out_activate_0_T_4 ? buffer_3_16 : _GEN_724; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_726 = 2'h3 == read_ptr[1:0] & 5'h11 == _io_out_activate_0_T_4 ? buffer_3_17 : _GEN_725; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_727 = 2'h3 == read_ptr[1:0] & 5'h12 == _io_out_activate_0_T_4 ? buffer_3_18 : _GEN_726; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_728 = 2'h3 == read_ptr[1:0] & 5'h13 == _io_out_activate_0_T_4 ? buffer_3_19 : _GEN_727; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_729 = 2'h3 == read_ptr[1:0] & 5'h14 == _io_out_activate_0_T_4 ? buffer_3_20 : _GEN_728; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_730 = 2'h3 == read_ptr[1:0] & 5'h15 == _io_out_activate_0_T_4 ? buffer_3_21 : _GEN_729; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_731 = 2'h3 == read_ptr[1:0] & 5'h16 == _io_out_activate_0_T_4 ? buffer_3_22 : _GEN_730; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_732 = 2'h3 == read_ptr[1:0] & 5'h17 == _io_out_activate_0_T_4 ? buffer_3_23 : _GEN_731; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_733 = 2'h3 == read_ptr[1:0] & 5'h18 == _io_out_activate_0_T_4 ? buffer_3_24 : _GEN_732; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_734 = 2'h3 == read_ptr[1:0] & 5'h19 == _io_out_activate_0_T_4 ? buffer_3_25 : _GEN_733; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_735 = 2'h3 == read_ptr[1:0] & 5'h1a == _io_out_activate_0_T_4 ? buffer_3_26 : _GEN_734; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_736 = 2'h3 == read_ptr[1:0] & 5'h1b == _io_out_activate_0_T_4 ? buffer_3_27 : _GEN_735; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_737 = 2'h3 == read_ptr[1:0] & 5'h1c == _io_out_activate_0_T_4 ? buffer_3_28 : _GEN_736; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_738 = 2'h3 == read_ptr[1:0] & 5'h1d == _io_out_activate_0_T_4 ? buffer_3_29 : _GEN_737; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_739 = 2'h3 == read_ptr[1:0] & 5'h1e == _io_out_activate_0_T_4 ? buffer_3_30 : _GEN_738; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_740 = 2'h3 == read_ptr[1:0] & 5'h1f == _io_out_activate_0_T_4 ? buffer_3_31 : _GEN_739; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_741 = 2'h3 == read_ptr[1:0] & 6'h20 == _GEN_2645 ? buffer_3_32 : _GEN_740; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_742 = 2'h3 == read_ptr[1:0] & 6'h21 == _GEN_2645 ? buffer_3_33 : _GEN_741; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_743 = 2'h3 == read_ptr[1:0] & 6'h22 == _GEN_2645 ? buffer_3_34 : _GEN_742; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_744 = 2'h3 == read_ptr[1:0] & 6'h23 == _GEN_2645 ? buffer_3_35 : _GEN_743; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_745 = 2'h3 == read_ptr[1:0] & 6'h24 == _GEN_2645 ? buffer_3_36 : _GEN_744; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_746 = 2'h3 == read_ptr[1:0] & 6'h25 == _GEN_2645 ? buffer_3_37 : _GEN_745; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_747 = 2'h3 == read_ptr[1:0] & 6'h26 == _GEN_2645 ? buffer_3_38 : _GEN_746; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_748 = 2'h3 == read_ptr[1:0] & 6'h27 == _GEN_2645 ? buffer_3_39 : _GEN_747; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_749 = 2'h3 == read_ptr[1:0] & 6'h28 == _GEN_2645 ? buffer_3_40 : _GEN_748; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_750 = 2'h3 == read_ptr[1:0] & 6'h29 == _GEN_2645 ? buffer_3_41 : _GEN_749; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_751 = 2'h3 == read_ptr[1:0] & 6'h2a == _GEN_2645 ? buffer_3_42 : _GEN_750; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_752 = 2'h3 == read_ptr[1:0] & 6'h2b == _GEN_2645 ? buffer_3_43 : _GEN_751; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_753 = 2'h3 == read_ptr[1:0] & 6'h2c == _GEN_2645 ? buffer_3_44 : _GEN_752; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_754 = 2'h3 == read_ptr[1:0] & 6'h2d == _GEN_2645 ? buffer_3_45 : _GEN_753; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_755 = 2'h3 == read_ptr[1:0] & 6'h2e == _GEN_2645 ? buffer_3_46 : _GEN_754; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_756 = 2'h3 == read_ptr[1:0] & 6'h2f == _GEN_2645 ? buffer_3_47 : _GEN_755; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_757 = 2'h3 == read_ptr[1:0] & 6'h30 == _GEN_2645 ? buffer_3_48 : _GEN_756; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_758 = 2'h3 == read_ptr[1:0] & 6'h31 == _GEN_2645 ? buffer_3_49 : _GEN_757; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_759 = 2'h3 == read_ptr[1:0] & 6'h32 == _GEN_2645 ? buffer_3_50 : _GEN_758; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_760 = 2'h3 == read_ptr[1:0] & 6'h33 == _GEN_2645 ? buffer_3_51 : _GEN_759; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_761 = 2'h3 == read_ptr[1:0] & 6'h34 == _GEN_2645 ? buffer_3_52 : _GEN_760; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_762 = 2'h3 == read_ptr[1:0] & 6'h35 == _GEN_2645 ? buffer_3_53 : _GEN_761; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_763 = 2'h3 == read_ptr[1:0] & 6'h36 == _GEN_2645 ? buffer_3_54 : _GEN_762; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_764 = 2'h3 == read_ptr[1:0] & 6'h37 == _GEN_2645 ? buffer_3_55 : _GEN_763; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_765 = 2'h3 == read_ptr[1:0] & 6'h38 == _GEN_2645 ? buffer_3_56 : _GEN_764; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_766 = 2'h3 == read_ptr[1:0] & 6'h39 == _GEN_2645 ? buffer_3_57 : _GEN_765; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_767 = 2'h3 == read_ptr[1:0] & 6'h3a == _GEN_2645 ? buffer_3_58 : _GEN_766; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_768 = 2'h3 == read_ptr[1:0] & 6'h3b == _GEN_2645 ? buffer_3_59 : _GEN_767; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_769 = 2'h3 == read_ptr[1:0] & 6'h3c == _GEN_2645 ? buffer_3_60 : _GEN_768; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_770 = 2'h3 == read_ptr[1:0] & 6'h3d == _GEN_2645 ? buffer_3_61 : _GEN_769; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_771 = 2'h3 == read_ptr[1:0] & 6'h3e == _GEN_2645 ? buffer_3_62 : _GEN_770; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_772 = 2'h3 == read_ptr[1:0] & 6'h3f == _GEN_2645 ? buffer_3_63 : _GEN_771; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_773 = 5'h0 < flow_ptr & flow_ptr <= 5'h8 ? _GEN_772 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [4:0] _io_out_activate_1_T_2 = 5'h8 + flow_ptr; // @[Activation_Buffer.scala 76:88]
  wire [4:0] _io_out_activate_1_T_4 = _io_out_activate_1_T_2 - 5'h2; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_775 = 2'h0 == read_ptr[1:0] & 5'h1 == _io_out_activate_1_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_776 = 2'h0 == read_ptr[1:0] & 5'h2 == _io_out_activate_1_T_4 ? buffer_0_2 : _GEN_775; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_777 = 2'h0 == read_ptr[1:0] & 5'h3 == _io_out_activate_1_T_4 ? buffer_0_3 : _GEN_776; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_778 = 2'h0 == read_ptr[1:0] & 5'h4 == _io_out_activate_1_T_4 ? buffer_0_4 : _GEN_777; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_779 = 2'h0 == read_ptr[1:0] & 5'h5 == _io_out_activate_1_T_4 ? buffer_0_5 : _GEN_778; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_780 = 2'h0 == read_ptr[1:0] & 5'h6 == _io_out_activate_1_T_4 ? buffer_0_6 : _GEN_779; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_781 = 2'h0 == read_ptr[1:0] & 5'h7 == _io_out_activate_1_T_4 ? buffer_0_7 : _GEN_780; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_782 = 2'h0 == read_ptr[1:0] & 5'h8 == _io_out_activate_1_T_4 ? buffer_0_8 : _GEN_781; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_783 = 2'h0 == read_ptr[1:0] & 5'h9 == _io_out_activate_1_T_4 ? buffer_0_9 : _GEN_782; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_784 = 2'h0 == read_ptr[1:0] & 5'ha == _io_out_activate_1_T_4 ? buffer_0_10 : _GEN_783; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_785 = 2'h0 == read_ptr[1:0] & 5'hb == _io_out_activate_1_T_4 ? buffer_0_11 : _GEN_784; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_786 = 2'h0 == read_ptr[1:0] & 5'hc == _io_out_activate_1_T_4 ? buffer_0_12 : _GEN_785; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_787 = 2'h0 == read_ptr[1:0] & 5'hd == _io_out_activate_1_T_4 ? buffer_0_13 : _GEN_786; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_788 = 2'h0 == read_ptr[1:0] & 5'he == _io_out_activate_1_T_4 ? buffer_0_14 : _GEN_787; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_789 = 2'h0 == read_ptr[1:0] & 5'hf == _io_out_activate_1_T_4 ? buffer_0_15 : _GEN_788; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_790 = 2'h0 == read_ptr[1:0] & 5'h10 == _io_out_activate_1_T_4 ? buffer_0_16 : _GEN_789; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_791 = 2'h0 == read_ptr[1:0] & 5'h11 == _io_out_activate_1_T_4 ? buffer_0_17 : _GEN_790; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_792 = 2'h0 == read_ptr[1:0] & 5'h12 == _io_out_activate_1_T_4 ? buffer_0_18 : _GEN_791; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_793 = 2'h0 == read_ptr[1:0] & 5'h13 == _io_out_activate_1_T_4 ? buffer_0_19 : _GEN_792; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_794 = 2'h0 == read_ptr[1:0] & 5'h14 == _io_out_activate_1_T_4 ? buffer_0_20 : _GEN_793; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_795 = 2'h0 == read_ptr[1:0] & 5'h15 == _io_out_activate_1_T_4 ? buffer_0_21 : _GEN_794; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_796 = 2'h0 == read_ptr[1:0] & 5'h16 == _io_out_activate_1_T_4 ? buffer_0_22 : _GEN_795; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_797 = 2'h0 == read_ptr[1:0] & 5'h17 == _io_out_activate_1_T_4 ? buffer_0_23 : _GEN_796; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_798 = 2'h0 == read_ptr[1:0] & 5'h18 == _io_out_activate_1_T_4 ? buffer_0_24 : _GEN_797; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_799 = 2'h0 == read_ptr[1:0] & 5'h19 == _io_out_activate_1_T_4 ? buffer_0_25 : _GEN_798; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_800 = 2'h0 == read_ptr[1:0] & 5'h1a == _io_out_activate_1_T_4 ? buffer_0_26 : _GEN_799; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_801 = 2'h0 == read_ptr[1:0] & 5'h1b == _io_out_activate_1_T_4 ? buffer_0_27 : _GEN_800; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_802 = 2'h0 == read_ptr[1:0] & 5'h1c == _io_out_activate_1_T_4 ? buffer_0_28 : _GEN_801; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_803 = 2'h0 == read_ptr[1:0] & 5'h1d == _io_out_activate_1_T_4 ? buffer_0_29 : _GEN_802; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_804 = 2'h0 == read_ptr[1:0] & 5'h1e == _io_out_activate_1_T_4 ? buffer_0_30 : _GEN_803; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_805 = 2'h0 == read_ptr[1:0] & 5'h1f == _io_out_activate_1_T_4 ? buffer_0_31 : _GEN_804; // @[Activation_Buffer.scala 76:{28,28}]
  wire [5:0] _GEN_3283 = {{1'd0}, _io_out_activate_1_T_4}; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_806 = 2'h0 == read_ptr[1:0] & 6'h20 == _GEN_3283 ? buffer_0_32 : _GEN_805; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_807 = 2'h0 == read_ptr[1:0] & 6'h21 == _GEN_3283 ? buffer_0_33 : _GEN_806; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_808 = 2'h0 == read_ptr[1:0] & 6'h22 == _GEN_3283 ? buffer_0_34 : _GEN_807; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_809 = 2'h0 == read_ptr[1:0] & 6'h23 == _GEN_3283 ? buffer_0_35 : _GEN_808; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_810 = 2'h0 == read_ptr[1:0] & 6'h24 == _GEN_3283 ? buffer_0_36 : _GEN_809; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_811 = 2'h0 == read_ptr[1:0] & 6'h25 == _GEN_3283 ? buffer_0_37 : _GEN_810; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_812 = 2'h0 == read_ptr[1:0] & 6'h26 == _GEN_3283 ? buffer_0_38 : _GEN_811; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_813 = 2'h0 == read_ptr[1:0] & 6'h27 == _GEN_3283 ? buffer_0_39 : _GEN_812; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_814 = 2'h0 == read_ptr[1:0] & 6'h28 == _GEN_3283 ? buffer_0_40 : _GEN_813; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_815 = 2'h0 == read_ptr[1:0] & 6'h29 == _GEN_3283 ? buffer_0_41 : _GEN_814; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_816 = 2'h0 == read_ptr[1:0] & 6'h2a == _GEN_3283 ? buffer_0_42 : _GEN_815; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_817 = 2'h0 == read_ptr[1:0] & 6'h2b == _GEN_3283 ? buffer_0_43 : _GEN_816; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_818 = 2'h0 == read_ptr[1:0] & 6'h2c == _GEN_3283 ? buffer_0_44 : _GEN_817; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_819 = 2'h0 == read_ptr[1:0] & 6'h2d == _GEN_3283 ? buffer_0_45 : _GEN_818; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_820 = 2'h0 == read_ptr[1:0] & 6'h2e == _GEN_3283 ? buffer_0_46 : _GEN_819; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_821 = 2'h0 == read_ptr[1:0] & 6'h2f == _GEN_3283 ? buffer_0_47 : _GEN_820; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_822 = 2'h0 == read_ptr[1:0] & 6'h30 == _GEN_3283 ? buffer_0_48 : _GEN_821; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_823 = 2'h0 == read_ptr[1:0] & 6'h31 == _GEN_3283 ? buffer_0_49 : _GEN_822; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_824 = 2'h0 == read_ptr[1:0] & 6'h32 == _GEN_3283 ? buffer_0_50 : _GEN_823; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_825 = 2'h0 == read_ptr[1:0] & 6'h33 == _GEN_3283 ? buffer_0_51 : _GEN_824; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_826 = 2'h0 == read_ptr[1:0] & 6'h34 == _GEN_3283 ? buffer_0_52 : _GEN_825; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_827 = 2'h0 == read_ptr[1:0] & 6'h35 == _GEN_3283 ? buffer_0_53 : _GEN_826; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_828 = 2'h0 == read_ptr[1:0] & 6'h36 == _GEN_3283 ? buffer_0_54 : _GEN_827; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_829 = 2'h0 == read_ptr[1:0] & 6'h37 == _GEN_3283 ? buffer_0_55 : _GEN_828; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_830 = 2'h0 == read_ptr[1:0] & 6'h38 == _GEN_3283 ? buffer_0_56 : _GEN_829; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_831 = 2'h0 == read_ptr[1:0] & 6'h39 == _GEN_3283 ? buffer_0_57 : _GEN_830; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_832 = 2'h0 == read_ptr[1:0] & 6'h3a == _GEN_3283 ? buffer_0_58 : _GEN_831; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_833 = 2'h0 == read_ptr[1:0] & 6'h3b == _GEN_3283 ? buffer_0_59 : _GEN_832; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_834 = 2'h0 == read_ptr[1:0] & 6'h3c == _GEN_3283 ? buffer_0_60 : _GEN_833; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_835 = 2'h0 == read_ptr[1:0] & 6'h3d == _GEN_3283 ? buffer_0_61 : _GEN_834; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_836 = 2'h0 == read_ptr[1:0] & 6'h3e == _GEN_3283 ? buffer_0_62 : _GEN_835; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_837 = 2'h0 == read_ptr[1:0] & 6'h3f == _GEN_3283 ? buffer_0_63 : _GEN_836; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_838 = 2'h1 == read_ptr[1:0] & 5'h0 == _io_out_activate_1_T_4 ? buffer_1_0 : _GEN_837; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_839 = 2'h1 == read_ptr[1:0] & 5'h1 == _io_out_activate_1_T_4 ? buffer_1_1 : _GEN_838; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_840 = 2'h1 == read_ptr[1:0] & 5'h2 == _io_out_activate_1_T_4 ? buffer_1_2 : _GEN_839; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_841 = 2'h1 == read_ptr[1:0] & 5'h3 == _io_out_activate_1_T_4 ? buffer_1_3 : _GEN_840; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_842 = 2'h1 == read_ptr[1:0] & 5'h4 == _io_out_activate_1_T_4 ? buffer_1_4 : _GEN_841; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_843 = 2'h1 == read_ptr[1:0] & 5'h5 == _io_out_activate_1_T_4 ? buffer_1_5 : _GEN_842; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_844 = 2'h1 == read_ptr[1:0] & 5'h6 == _io_out_activate_1_T_4 ? buffer_1_6 : _GEN_843; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_845 = 2'h1 == read_ptr[1:0] & 5'h7 == _io_out_activate_1_T_4 ? buffer_1_7 : _GEN_844; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_846 = 2'h1 == read_ptr[1:0] & 5'h8 == _io_out_activate_1_T_4 ? buffer_1_8 : _GEN_845; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_847 = 2'h1 == read_ptr[1:0] & 5'h9 == _io_out_activate_1_T_4 ? buffer_1_9 : _GEN_846; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_848 = 2'h1 == read_ptr[1:0] & 5'ha == _io_out_activate_1_T_4 ? buffer_1_10 : _GEN_847; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_849 = 2'h1 == read_ptr[1:0] & 5'hb == _io_out_activate_1_T_4 ? buffer_1_11 : _GEN_848; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_850 = 2'h1 == read_ptr[1:0] & 5'hc == _io_out_activate_1_T_4 ? buffer_1_12 : _GEN_849; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_851 = 2'h1 == read_ptr[1:0] & 5'hd == _io_out_activate_1_T_4 ? buffer_1_13 : _GEN_850; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_852 = 2'h1 == read_ptr[1:0] & 5'he == _io_out_activate_1_T_4 ? buffer_1_14 : _GEN_851; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_853 = 2'h1 == read_ptr[1:0] & 5'hf == _io_out_activate_1_T_4 ? buffer_1_15 : _GEN_852; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_854 = 2'h1 == read_ptr[1:0] & 5'h10 == _io_out_activate_1_T_4 ? buffer_1_16 : _GEN_853; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_855 = 2'h1 == read_ptr[1:0] & 5'h11 == _io_out_activate_1_T_4 ? buffer_1_17 : _GEN_854; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_856 = 2'h1 == read_ptr[1:0] & 5'h12 == _io_out_activate_1_T_4 ? buffer_1_18 : _GEN_855; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_857 = 2'h1 == read_ptr[1:0] & 5'h13 == _io_out_activate_1_T_4 ? buffer_1_19 : _GEN_856; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_858 = 2'h1 == read_ptr[1:0] & 5'h14 == _io_out_activate_1_T_4 ? buffer_1_20 : _GEN_857; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_859 = 2'h1 == read_ptr[1:0] & 5'h15 == _io_out_activate_1_T_4 ? buffer_1_21 : _GEN_858; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_860 = 2'h1 == read_ptr[1:0] & 5'h16 == _io_out_activate_1_T_4 ? buffer_1_22 : _GEN_859; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_861 = 2'h1 == read_ptr[1:0] & 5'h17 == _io_out_activate_1_T_4 ? buffer_1_23 : _GEN_860; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_862 = 2'h1 == read_ptr[1:0] & 5'h18 == _io_out_activate_1_T_4 ? buffer_1_24 : _GEN_861; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_863 = 2'h1 == read_ptr[1:0] & 5'h19 == _io_out_activate_1_T_4 ? buffer_1_25 : _GEN_862; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_864 = 2'h1 == read_ptr[1:0] & 5'h1a == _io_out_activate_1_T_4 ? buffer_1_26 : _GEN_863; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_865 = 2'h1 == read_ptr[1:0] & 5'h1b == _io_out_activate_1_T_4 ? buffer_1_27 : _GEN_864; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_866 = 2'h1 == read_ptr[1:0] & 5'h1c == _io_out_activate_1_T_4 ? buffer_1_28 : _GEN_865; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_867 = 2'h1 == read_ptr[1:0] & 5'h1d == _io_out_activate_1_T_4 ? buffer_1_29 : _GEN_866; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_868 = 2'h1 == read_ptr[1:0] & 5'h1e == _io_out_activate_1_T_4 ? buffer_1_30 : _GEN_867; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_869 = 2'h1 == read_ptr[1:0] & 5'h1f == _io_out_activate_1_T_4 ? buffer_1_31 : _GEN_868; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_870 = 2'h1 == read_ptr[1:0] & 6'h20 == _GEN_3283 ? buffer_1_32 : _GEN_869; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_871 = 2'h1 == read_ptr[1:0] & 6'h21 == _GEN_3283 ? buffer_1_33 : _GEN_870; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_872 = 2'h1 == read_ptr[1:0] & 6'h22 == _GEN_3283 ? buffer_1_34 : _GEN_871; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_873 = 2'h1 == read_ptr[1:0] & 6'h23 == _GEN_3283 ? buffer_1_35 : _GEN_872; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_874 = 2'h1 == read_ptr[1:0] & 6'h24 == _GEN_3283 ? buffer_1_36 : _GEN_873; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_875 = 2'h1 == read_ptr[1:0] & 6'h25 == _GEN_3283 ? buffer_1_37 : _GEN_874; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_876 = 2'h1 == read_ptr[1:0] & 6'h26 == _GEN_3283 ? buffer_1_38 : _GEN_875; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_877 = 2'h1 == read_ptr[1:0] & 6'h27 == _GEN_3283 ? buffer_1_39 : _GEN_876; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_878 = 2'h1 == read_ptr[1:0] & 6'h28 == _GEN_3283 ? buffer_1_40 : _GEN_877; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_879 = 2'h1 == read_ptr[1:0] & 6'h29 == _GEN_3283 ? buffer_1_41 : _GEN_878; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_880 = 2'h1 == read_ptr[1:0] & 6'h2a == _GEN_3283 ? buffer_1_42 : _GEN_879; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_881 = 2'h1 == read_ptr[1:0] & 6'h2b == _GEN_3283 ? buffer_1_43 : _GEN_880; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_882 = 2'h1 == read_ptr[1:0] & 6'h2c == _GEN_3283 ? buffer_1_44 : _GEN_881; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_883 = 2'h1 == read_ptr[1:0] & 6'h2d == _GEN_3283 ? buffer_1_45 : _GEN_882; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_884 = 2'h1 == read_ptr[1:0] & 6'h2e == _GEN_3283 ? buffer_1_46 : _GEN_883; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_885 = 2'h1 == read_ptr[1:0] & 6'h2f == _GEN_3283 ? buffer_1_47 : _GEN_884; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_886 = 2'h1 == read_ptr[1:0] & 6'h30 == _GEN_3283 ? buffer_1_48 : _GEN_885; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_887 = 2'h1 == read_ptr[1:0] & 6'h31 == _GEN_3283 ? buffer_1_49 : _GEN_886; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_888 = 2'h1 == read_ptr[1:0] & 6'h32 == _GEN_3283 ? buffer_1_50 : _GEN_887; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_889 = 2'h1 == read_ptr[1:0] & 6'h33 == _GEN_3283 ? buffer_1_51 : _GEN_888; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_890 = 2'h1 == read_ptr[1:0] & 6'h34 == _GEN_3283 ? buffer_1_52 : _GEN_889; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_891 = 2'h1 == read_ptr[1:0] & 6'h35 == _GEN_3283 ? buffer_1_53 : _GEN_890; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_892 = 2'h1 == read_ptr[1:0] & 6'h36 == _GEN_3283 ? buffer_1_54 : _GEN_891; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_893 = 2'h1 == read_ptr[1:0] & 6'h37 == _GEN_3283 ? buffer_1_55 : _GEN_892; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_894 = 2'h1 == read_ptr[1:0] & 6'h38 == _GEN_3283 ? buffer_1_56 : _GEN_893; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_895 = 2'h1 == read_ptr[1:0] & 6'h39 == _GEN_3283 ? buffer_1_57 : _GEN_894; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_896 = 2'h1 == read_ptr[1:0] & 6'h3a == _GEN_3283 ? buffer_1_58 : _GEN_895; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_897 = 2'h1 == read_ptr[1:0] & 6'h3b == _GEN_3283 ? buffer_1_59 : _GEN_896; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_898 = 2'h1 == read_ptr[1:0] & 6'h3c == _GEN_3283 ? buffer_1_60 : _GEN_897; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_899 = 2'h1 == read_ptr[1:0] & 6'h3d == _GEN_3283 ? buffer_1_61 : _GEN_898; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_900 = 2'h1 == read_ptr[1:0] & 6'h3e == _GEN_3283 ? buffer_1_62 : _GEN_899; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_901 = 2'h1 == read_ptr[1:0] & 6'h3f == _GEN_3283 ? buffer_1_63 : _GEN_900; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_902 = 2'h2 == read_ptr[1:0] & 5'h0 == _io_out_activate_1_T_4 ? buffer_2_0 : _GEN_901; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_903 = 2'h2 == read_ptr[1:0] & 5'h1 == _io_out_activate_1_T_4 ? buffer_2_1 : _GEN_902; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_904 = 2'h2 == read_ptr[1:0] & 5'h2 == _io_out_activate_1_T_4 ? buffer_2_2 : _GEN_903; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_905 = 2'h2 == read_ptr[1:0] & 5'h3 == _io_out_activate_1_T_4 ? buffer_2_3 : _GEN_904; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_906 = 2'h2 == read_ptr[1:0] & 5'h4 == _io_out_activate_1_T_4 ? buffer_2_4 : _GEN_905; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_907 = 2'h2 == read_ptr[1:0] & 5'h5 == _io_out_activate_1_T_4 ? buffer_2_5 : _GEN_906; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_908 = 2'h2 == read_ptr[1:0] & 5'h6 == _io_out_activate_1_T_4 ? buffer_2_6 : _GEN_907; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_909 = 2'h2 == read_ptr[1:0] & 5'h7 == _io_out_activate_1_T_4 ? buffer_2_7 : _GEN_908; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_910 = 2'h2 == read_ptr[1:0] & 5'h8 == _io_out_activate_1_T_4 ? buffer_2_8 : _GEN_909; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_911 = 2'h2 == read_ptr[1:0] & 5'h9 == _io_out_activate_1_T_4 ? buffer_2_9 : _GEN_910; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_912 = 2'h2 == read_ptr[1:0] & 5'ha == _io_out_activate_1_T_4 ? buffer_2_10 : _GEN_911; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_913 = 2'h2 == read_ptr[1:0] & 5'hb == _io_out_activate_1_T_4 ? buffer_2_11 : _GEN_912; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_914 = 2'h2 == read_ptr[1:0] & 5'hc == _io_out_activate_1_T_4 ? buffer_2_12 : _GEN_913; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_915 = 2'h2 == read_ptr[1:0] & 5'hd == _io_out_activate_1_T_4 ? buffer_2_13 : _GEN_914; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_916 = 2'h2 == read_ptr[1:0] & 5'he == _io_out_activate_1_T_4 ? buffer_2_14 : _GEN_915; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_917 = 2'h2 == read_ptr[1:0] & 5'hf == _io_out_activate_1_T_4 ? buffer_2_15 : _GEN_916; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_918 = 2'h2 == read_ptr[1:0] & 5'h10 == _io_out_activate_1_T_4 ? buffer_2_16 : _GEN_917; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_919 = 2'h2 == read_ptr[1:0] & 5'h11 == _io_out_activate_1_T_4 ? buffer_2_17 : _GEN_918; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_920 = 2'h2 == read_ptr[1:0] & 5'h12 == _io_out_activate_1_T_4 ? buffer_2_18 : _GEN_919; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_921 = 2'h2 == read_ptr[1:0] & 5'h13 == _io_out_activate_1_T_4 ? buffer_2_19 : _GEN_920; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_922 = 2'h2 == read_ptr[1:0] & 5'h14 == _io_out_activate_1_T_4 ? buffer_2_20 : _GEN_921; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_923 = 2'h2 == read_ptr[1:0] & 5'h15 == _io_out_activate_1_T_4 ? buffer_2_21 : _GEN_922; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_924 = 2'h2 == read_ptr[1:0] & 5'h16 == _io_out_activate_1_T_4 ? buffer_2_22 : _GEN_923; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_925 = 2'h2 == read_ptr[1:0] & 5'h17 == _io_out_activate_1_T_4 ? buffer_2_23 : _GEN_924; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_926 = 2'h2 == read_ptr[1:0] & 5'h18 == _io_out_activate_1_T_4 ? buffer_2_24 : _GEN_925; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_927 = 2'h2 == read_ptr[1:0] & 5'h19 == _io_out_activate_1_T_4 ? buffer_2_25 : _GEN_926; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_928 = 2'h2 == read_ptr[1:0] & 5'h1a == _io_out_activate_1_T_4 ? buffer_2_26 : _GEN_927; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_929 = 2'h2 == read_ptr[1:0] & 5'h1b == _io_out_activate_1_T_4 ? buffer_2_27 : _GEN_928; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_930 = 2'h2 == read_ptr[1:0] & 5'h1c == _io_out_activate_1_T_4 ? buffer_2_28 : _GEN_929; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_931 = 2'h2 == read_ptr[1:0] & 5'h1d == _io_out_activate_1_T_4 ? buffer_2_29 : _GEN_930; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_932 = 2'h2 == read_ptr[1:0] & 5'h1e == _io_out_activate_1_T_4 ? buffer_2_30 : _GEN_931; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_933 = 2'h2 == read_ptr[1:0] & 5'h1f == _io_out_activate_1_T_4 ? buffer_2_31 : _GEN_932; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_934 = 2'h2 == read_ptr[1:0] & 6'h20 == _GEN_3283 ? buffer_2_32 : _GEN_933; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_935 = 2'h2 == read_ptr[1:0] & 6'h21 == _GEN_3283 ? buffer_2_33 : _GEN_934; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_936 = 2'h2 == read_ptr[1:0] & 6'h22 == _GEN_3283 ? buffer_2_34 : _GEN_935; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_937 = 2'h2 == read_ptr[1:0] & 6'h23 == _GEN_3283 ? buffer_2_35 : _GEN_936; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_938 = 2'h2 == read_ptr[1:0] & 6'h24 == _GEN_3283 ? buffer_2_36 : _GEN_937; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_939 = 2'h2 == read_ptr[1:0] & 6'h25 == _GEN_3283 ? buffer_2_37 : _GEN_938; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_940 = 2'h2 == read_ptr[1:0] & 6'h26 == _GEN_3283 ? buffer_2_38 : _GEN_939; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_941 = 2'h2 == read_ptr[1:0] & 6'h27 == _GEN_3283 ? buffer_2_39 : _GEN_940; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_942 = 2'h2 == read_ptr[1:0] & 6'h28 == _GEN_3283 ? buffer_2_40 : _GEN_941; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_943 = 2'h2 == read_ptr[1:0] & 6'h29 == _GEN_3283 ? buffer_2_41 : _GEN_942; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_944 = 2'h2 == read_ptr[1:0] & 6'h2a == _GEN_3283 ? buffer_2_42 : _GEN_943; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_945 = 2'h2 == read_ptr[1:0] & 6'h2b == _GEN_3283 ? buffer_2_43 : _GEN_944; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_946 = 2'h2 == read_ptr[1:0] & 6'h2c == _GEN_3283 ? buffer_2_44 : _GEN_945; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_947 = 2'h2 == read_ptr[1:0] & 6'h2d == _GEN_3283 ? buffer_2_45 : _GEN_946; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_948 = 2'h2 == read_ptr[1:0] & 6'h2e == _GEN_3283 ? buffer_2_46 : _GEN_947; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_949 = 2'h2 == read_ptr[1:0] & 6'h2f == _GEN_3283 ? buffer_2_47 : _GEN_948; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_950 = 2'h2 == read_ptr[1:0] & 6'h30 == _GEN_3283 ? buffer_2_48 : _GEN_949; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_951 = 2'h2 == read_ptr[1:0] & 6'h31 == _GEN_3283 ? buffer_2_49 : _GEN_950; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_952 = 2'h2 == read_ptr[1:0] & 6'h32 == _GEN_3283 ? buffer_2_50 : _GEN_951; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_953 = 2'h2 == read_ptr[1:0] & 6'h33 == _GEN_3283 ? buffer_2_51 : _GEN_952; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_954 = 2'h2 == read_ptr[1:0] & 6'h34 == _GEN_3283 ? buffer_2_52 : _GEN_953; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_955 = 2'h2 == read_ptr[1:0] & 6'h35 == _GEN_3283 ? buffer_2_53 : _GEN_954; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_956 = 2'h2 == read_ptr[1:0] & 6'h36 == _GEN_3283 ? buffer_2_54 : _GEN_955; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_957 = 2'h2 == read_ptr[1:0] & 6'h37 == _GEN_3283 ? buffer_2_55 : _GEN_956; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_958 = 2'h2 == read_ptr[1:0] & 6'h38 == _GEN_3283 ? buffer_2_56 : _GEN_957; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_959 = 2'h2 == read_ptr[1:0] & 6'h39 == _GEN_3283 ? buffer_2_57 : _GEN_958; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_960 = 2'h2 == read_ptr[1:0] & 6'h3a == _GEN_3283 ? buffer_2_58 : _GEN_959; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_961 = 2'h2 == read_ptr[1:0] & 6'h3b == _GEN_3283 ? buffer_2_59 : _GEN_960; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_962 = 2'h2 == read_ptr[1:0] & 6'h3c == _GEN_3283 ? buffer_2_60 : _GEN_961; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_963 = 2'h2 == read_ptr[1:0] & 6'h3d == _GEN_3283 ? buffer_2_61 : _GEN_962; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_964 = 2'h2 == read_ptr[1:0] & 6'h3e == _GEN_3283 ? buffer_2_62 : _GEN_963; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_965 = 2'h2 == read_ptr[1:0] & 6'h3f == _GEN_3283 ? buffer_2_63 : _GEN_964; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_966 = 2'h3 == read_ptr[1:0] & 5'h0 == _io_out_activate_1_T_4 ? buffer_3_0 : _GEN_965; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_967 = 2'h3 == read_ptr[1:0] & 5'h1 == _io_out_activate_1_T_4 ? buffer_3_1 : _GEN_966; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_968 = 2'h3 == read_ptr[1:0] & 5'h2 == _io_out_activate_1_T_4 ? buffer_3_2 : _GEN_967; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_969 = 2'h3 == read_ptr[1:0] & 5'h3 == _io_out_activate_1_T_4 ? buffer_3_3 : _GEN_968; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_970 = 2'h3 == read_ptr[1:0] & 5'h4 == _io_out_activate_1_T_4 ? buffer_3_4 : _GEN_969; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_971 = 2'h3 == read_ptr[1:0] & 5'h5 == _io_out_activate_1_T_4 ? buffer_3_5 : _GEN_970; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_972 = 2'h3 == read_ptr[1:0] & 5'h6 == _io_out_activate_1_T_4 ? buffer_3_6 : _GEN_971; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_973 = 2'h3 == read_ptr[1:0] & 5'h7 == _io_out_activate_1_T_4 ? buffer_3_7 : _GEN_972; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_974 = 2'h3 == read_ptr[1:0] & 5'h8 == _io_out_activate_1_T_4 ? buffer_3_8 : _GEN_973; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_975 = 2'h3 == read_ptr[1:0] & 5'h9 == _io_out_activate_1_T_4 ? buffer_3_9 : _GEN_974; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_976 = 2'h3 == read_ptr[1:0] & 5'ha == _io_out_activate_1_T_4 ? buffer_3_10 : _GEN_975; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_977 = 2'h3 == read_ptr[1:0] & 5'hb == _io_out_activate_1_T_4 ? buffer_3_11 : _GEN_976; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_978 = 2'h3 == read_ptr[1:0] & 5'hc == _io_out_activate_1_T_4 ? buffer_3_12 : _GEN_977; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_979 = 2'h3 == read_ptr[1:0] & 5'hd == _io_out_activate_1_T_4 ? buffer_3_13 : _GEN_978; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_980 = 2'h3 == read_ptr[1:0] & 5'he == _io_out_activate_1_T_4 ? buffer_3_14 : _GEN_979; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_981 = 2'h3 == read_ptr[1:0] & 5'hf == _io_out_activate_1_T_4 ? buffer_3_15 : _GEN_980; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_982 = 2'h3 == read_ptr[1:0] & 5'h10 == _io_out_activate_1_T_4 ? buffer_3_16 : _GEN_981; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_983 = 2'h3 == read_ptr[1:0] & 5'h11 == _io_out_activate_1_T_4 ? buffer_3_17 : _GEN_982; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_984 = 2'h3 == read_ptr[1:0] & 5'h12 == _io_out_activate_1_T_4 ? buffer_3_18 : _GEN_983; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_985 = 2'h3 == read_ptr[1:0] & 5'h13 == _io_out_activate_1_T_4 ? buffer_3_19 : _GEN_984; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_986 = 2'h3 == read_ptr[1:0] & 5'h14 == _io_out_activate_1_T_4 ? buffer_3_20 : _GEN_985; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_987 = 2'h3 == read_ptr[1:0] & 5'h15 == _io_out_activate_1_T_4 ? buffer_3_21 : _GEN_986; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_988 = 2'h3 == read_ptr[1:0] & 5'h16 == _io_out_activate_1_T_4 ? buffer_3_22 : _GEN_987; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_989 = 2'h3 == read_ptr[1:0] & 5'h17 == _io_out_activate_1_T_4 ? buffer_3_23 : _GEN_988; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_990 = 2'h3 == read_ptr[1:0] & 5'h18 == _io_out_activate_1_T_4 ? buffer_3_24 : _GEN_989; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_991 = 2'h3 == read_ptr[1:0] & 5'h19 == _io_out_activate_1_T_4 ? buffer_3_25 : _GEN_990; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_992 = 2'h3 == read_ptr[1:0] & 5'h1a == _io_out_activate_1_T_4 ? buffer_3_26 : _GEN_991; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_993 = 2'h3 == read_ptr[1:0] & 5'h1b == _io_out_activate_1_T_4 ? buffer_3_27 : _GEN_992; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_994 = 2'h3 == read_ptr[1:0] & 5'h1c == _io_out_activate_1_T_4 ? buffer_3_28 : _GEN_993; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_995 = 2'h3 == read_ptr[1:0] & 5'h1d == _io_out_activate_1_T_4 ? buffer_3_29 : _GEN_994; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_996 = 2'h3 == read_ptr[1:0] & 5'h1e == _io_out_activate_1_T_4 ? buffer_3_30 : _GEN_995; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_997 = 2'h3 == read_ptr[1:0] & 5'h1f == _io_out_activate_1_T_4 ? buffer_3_31 : _GEN_996; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_998 = 2'h3 == read_ptr[1:0] & 6'h20 == _GEN_3283 ? buffer_3_32 : _GEN_997; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_999 = 2'h3 == read_ptr[1:0] & 6'h21 == _GEN_3283 ? buffer_3_33 : _GEN_998; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1000 = 2'h3 == read_ptr[1:0] & 6'h22 == _GEN_3283 ? buffer_3_34 : _GEN_999; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1001 = 2'h3 == read_ptr[1:0] & 6'h23 == _GEN_3283 ? buffer_3_35 : _GEN_1000; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1002 = 2'h3 == read_ptr[1:0] & 6'h24 == _GEN_3283 ? buffer_3_36 : _GEN_1001; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1003 = 2'h3 == read_ptr[1:0] & 6'h25 == _GEN_3283 ? buffer_3_37 : _GEN_1002; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1004 = 2'h3 == read_ptr[1:0] & 6'h26 == _GEN_3283 ? buffer_3_38 : _GEN_1003; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1005 = 2'h3 == read_ptr[1:0] & 6'h27 == _GEN_3283 ? buffer_3_39 : _GEN_1004; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1006 = 2'h3 == read_ptr[1:0] & 6'h28 == _GEN_3283 ? buffer_3_40 : _GEN_1005; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1007 = 2'h3 == read_ptr[1:0] & 6'h29 == _GEN_3283 ? buffer_3_41 : _GEN_1006; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1008 = 2'h3 == read_ptr[1:0] & 6'h2a == _GEN_3283 ? buffer_3_42 : _GEN_1007; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1009 = 2'h3 == read_ptr[1:0] & 6'h2b == _GEN_3283 ? buffer_3_43 : _GEN_1008; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1010 = 2'h3 == read_ptr[1:0] & 6'h2c == _GEN_3283 ? buffer_3_44 : _GEN_1009; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1011 = 2'h3 == read_ptr[1:0] & 6'h2d == _GEN_3283 ? buffer_3_45 : _GEN_1010; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1012 = 2'h3 == read_ptr[1:0] & 6'h2e == _GEN_3283 ? buffer_3_46 : _GEN_1011; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1013 = 2'h3 == read_ptr[1:0] & 6'h2f == _GEN_3283 ? buffer_3_47 : _GEN_1012; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1014 = 2'h3 == read_ptr[1:0] & 6'h30 == _GEN_3283 ? buffer_3_48 : _GEN_1013; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1015 = 2'h3 == read_ptr[1:0] & 6'h31 == _GEN_3283 ? buffer_3_49 : _GEN_1014; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1016 = 2'h3 == read_ptr[1:0] & 6'h32 == _GEN_3283 ? buffer_3_50 : _GEN_1015; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1017 = 2'h3 == read_ptr[1:0] & 6'h33 == _GEN_3283 ? buffer_3_51 : _GEN_1016; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1018 = 2'h3 == read_ptr[1:0] & 6'h34 == _GEN_3283 ? buffer_3_52 : _GEN_1017; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1019 = 2'h3 == read_ptr[1:0] & 6'h35 == _GEN_3283 ? buffer_3_53 : _GEN_1018; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1020 = 2'h3 == read_ptr[1:0] & 6'h36 == _GEN_3283 ? buffer_3_54 : _GEN_1019; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1021 = 2'h3 == read_ptr[1:0] & 6'h37 == _GEN_3283 ? buffer_3_55 : _GEN_1020; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1022 = 2'h3 == read_ptr[1:0] & 6'h38 == _GEN_3283 ? buffer_3_56 : _GEN_1021; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1023 = 2'h3 == read_ptr[1:0] & 6'h39 == _GEN_3283 ? buffer_3_57 : _GEN_1022; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1024 = 2'h3 == read_ptr[1:0] & 6'h3a == _GEN_3283 ? buffer_3_58 : _GEN_1023; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1025 = 2'h3 == read_ptr[1:0] & 6'h3b == _GEN_3283 ? buffer_3_59 : _GEN_1024; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1026 = 2'h3 == read_ptr[1:0] & 6'h3c == _GEN_3283 ? buffer_3_60 : _GEN_1025; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1027 = 2'h3 == read_ptr[1:0] & 6'h3d == _GEN_3283 ? buffer_3_61 : _GEN_1026; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1028 = 2'h3 == read_ptr[1:0] & 6'h3e == _GEN_3283 ? buffer_3_62 : _GEN_1027; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1029 = 2'h3 == read_ptr[1:0] & 6'h3f == _GEN_3283 ? buffer_3_63 : _GEN_1028; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1030 = 5'h1 < flow_ptr & flow_ptr <= 5'h9 ? _GEN_1029 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [4:0] _io_out_activate_2_T_2 = 5'h10 + flow_ptr; // @[Activation_Buffer.scala 76:88]
  wire [4:0] _io_out_activate_2_T_4 = _io_out_activate_2_T_2 - 5'h3; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_1032 = 2'h0 == read_ptr[1:0] & 5'h1 == _io_out_activate_2_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1033 = 2'h0 == read_ptr[1:0] & 5'h2 == _io_out_activate_2_T_4 ? buffer_0_2 : _GEN_1032; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1034 = 2'h0 == read_ptr[1:0] & 5'h3 == _io_out_activate_2_T_4 ? buffer_0_3 : _GEN_1033; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1035 = 2'h0 == read_ptr[1:0] & 5'h4 == _io_out_activate_2_T_4 ? buffer_0_4 : _GEN_1034; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1036 = 2'h0 == read_ptr[1:0] & 5'h5 == _io_out_activate_2_T_4 ? buffer_0_5 : _GEN_1035; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1037 = 2'h0 == read_ptr[1:0] & 5'h6 == _io_out_activate_2_T_4 ? buffer_0_6 : _GEN_1036; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1038 = 2'h0 == read_ptr[1:0] & 5'h7 == _io_out_activate_2_T_4 ? buffer_0_7 : _GEN_1037; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1039 = 2'h0 == read_ptr[1:0] & 5'h8 == _io_out_activate_2_T_4 ? buffer_0_8 : _GEN_1038; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1040 = 2'h0 == read_ptr[1:0] & 5'h9 == _io_out_activate_2_T_4 ? buffer_0_9 : _GEN_1039; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1041 = 2'h0 == read_ptr[1:0] & 5'ha == _io_out_activate_2_T_4 ? buffer_0_10 : _GEN_1040; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1042 = 2'h0 == read_ptr[1:0] & 5'hb == _io_out_activate_2_T_4 ? buffer_0_11 : _GEN_1041; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1043 = 2'h0 == read_ptr[1:0] & 5'hc == _io_out_activate_2_T_4 ? buffer_0_12 : _GEN_1042; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1044 = 2'h0 == read_ptr[1:0] & 5'hd == _io_out_activate_2_T_4 ? buffer_0_13 : _GEN_1043; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1045 = 2'h0 == read_ptr[1:0] & 5'he == _io_out_activate_2_T_4 ? buffer_0_14 : _GEN_1044; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1046 = 2'h0 == read_ptr[1:0] & 5'hf == _io_out_activate_2_T_4 ? buffer_0_15 : _GEN_1045; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1047 = 2'h0 == read_ptr[1:0] & 5'h10 == _io_out_activate_2_T_4 ? buffer_0_16 : _GEN_1046; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1048 = 2'h0 == read_ptr[1:0] & 5'h11 == _io_out_activate_2_T_4 ? buffer_0_17 : _GEN_1047; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1049 = 2'h0 == read_ptr[1:0] & 5'h12 == _io_out_activate_2_T_4 ? buffer_0_18 : _GEN_1048; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1050 = 2'h0 == read_ptr[1:0] & 5'h13 == _io_out_activate_2_T_4 ? buffer_0_19 : _GEN_1049; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1051 = 2'h0 == read_ptr[1:0] & 5'h14 == _io_out_activate_2_T_4 ? buffer_0_20 : _GEN_1050; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1052 = 2'h0 == read_ptr[1:0] & 5'h15 == _io_out_activate_2_T_4 ? buffer_0_21 : _GEN_1051; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1053 = 2'h0 == read_ptr[1:0] & 5'h16 == _io_out_activate_2_T_4 ? buffer_0_22 : _GEN_1052; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1054 = 2'h0 == read_ptr[1:0] & 5'h17 == _io_out_activate_2_T_4 ? buffer_0_23 : _GEN_1053; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1055 = 2'h0 == read_ptr[1:0] & 5'h18 == _io_out_activate_2_T_4 ? buffer_0_24 : _GEN_1054; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1056 = 2'h0 == read_ptr[1:0] & 5'h19 == _io_out_activate_2_T_4 ? buffer_0_25 : _GEN_1055; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1057 = 2'h0 == read_ptr[1:0] & 5'h1a == _io_out_activate_2_T_4 ? buffer_0_26 : _GEN_1056; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1058 = 2'h0 == read_ptr[1:0] & 5'h1b == _io_out_activate_2_T_4 ? buffer_0_27 : _GEN_1057; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1059 = 2'h0 == read_ptr[1:0] & 5'h1c == _io_out_activate_2_T_4 ? buffer_0_28 : _GEN_1058; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1060 = 2'h0 == read_ptr[1:0] & 5'h1d == _io_out_activate_2_T_4 ? buffer_0_29 : _GEN_1059; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1061 = 2'h0 == read_ptr[1:0] & 5'h1e == _io_out_activate_2_T_4 ? buffer_0_30 : _GEN_1060; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1062 = 2'h0 == read_ptr[1:0] & 5'h1f == _io_out_activate_2_T_4 ? buffer_0_31 : _GEN_1061; // @[Activation_Buffer.scala 76:{28,28}]
  wire [5:0] _GEN_3921 = {{1'd0}, _io_out_activate_2_T_4}; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1063 = 2'h0 == read_ptr[1:0] & 6'h20 == _GEN_3921 ? buffer_0_32 : _GEN_1062; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1064 = 2'h0 == read_ptr[1:0] & 6'h21 == _GEN_3921 ? buffer_0_33 : _GEN_1063; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1065 = 2'h0 == read_ptr[1:0] & 6'h22 == _GEN_3921 ? buffer_0_34 : _GEN_1064; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1066 = 2'h0 == read_ptr[1:0] & 6'h23 == _GEN_3921 ? buffer_0_35 : _GEN_1065; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1067 = 2'h0 == read_ptr[1:0] & 6'h24 == _GEN_3921 ? buffer_0_36 : _GEN_1066; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1068 = 2'h0 == read_ptr[1:0] & 6'h25 == _GEN_3921 ? buffer_0_37 : _GEN_1067; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1069 = 2'h0 == read_ptr[1:0] & 6'h26 == _GEN_3921 ? buffer_0_38 : _GEN_1068; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1070 = 2'h0 == read_ptr[1:0] & 6'h27 == _GEN_3921 ? buffer_0_39 : _GEN_1069; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1071 = 2'h0 == read_ptr[1:0] & 6'h28 == _GEN_3921 ? buffer_0_40 : _GEN_1070; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1072 = 2'h0 == read_ptr[1:0] & 6'h29 == _GEN_3921 ? buffer_0_41 : _GEN_1071; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1073 = 2'h0 == read_ptr[1:0] & 6'h2a == _GEN_3921 ? buffer_0_42 : _GEN_1072; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1074 = 2'h0 == read_ptr[1:0] & 6'h2b == _GEN_3921 ? buffer_0_43 : _GEN_1073; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1075 = 2'h0 == read_ptr[1:0] & 6'h2c == _GEN_3921 ? buffer_0_44 : _GEN_1074; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1076 = 2'h0 == read_ptr[1:0] & 6'h2d == _GEN_3921 ? buffer_0_45 : _GEN_1075; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1077 = 2'h0 == read_ptr[1:0] & 6'h2e == _GEN_3921 ? buffer_0_46 : _GEN_1076; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1078 = 2'h0 == read_ptr[1:0] & 6'h2f == _GEN_3921 ? buffer_0_47 : _GEN_1077; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1079 = 2'h0 == read_ptr[1:0] & 6'h30 == _GEN_3921 ? buffer_0_48 : _GEN_1078; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1080 = 2'h0 == read_ptr[1:0] & 6'h31 == _GEN_3921 ? buffer_0_49 : _GEN_1079; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1081 = 2'h0 == read_ptr[1:0] & 6'h32 == _GEN_3921 ? buffer_0_50 : _GEN_1080; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1082 = 2'h0 == read_ptr[1:0] & 6'h33 == _GEN_3921 ? buffer_0_51 : _GEN_1081; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1083 = 2'h0 == read_ptr[1:0] & 6'h34 == _GEN_3921 ? buffer_0_52 : _GEN_1082; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1084 = 2'h0 == read_ptr[1:0] & 6'h35 == _GEN_3921 ? buffer_0_53 : _GEN_1083; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1085 = 2'h0 == read_ptr[1:0] & 6'h36 == _GEN_3921 ? buffer_0_54 : _GEN_1084; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1086 = 2'h0 == read_ptr[1:0] & 6'h37 == _GEN_3921 ? buffer_0_55 : _GEN_1085; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1087 = 2'h0 == read_ptr[1:0] & 6'h38 == _GEN_3921 ? buffer_0_56 : _GEN_1086; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1088 = 2'h0 == read_ptr[1:0] & 6'h39 == _GEN_3921 ? buffer_0_57 : _GEN_1087; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1089 = 2'h0 == read_ptr[1:0] & 6'h3a == _GEN_3921 ? buffer_0_58 : _GEN_1088; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1090 = 2'h0 == read_ptr[1:0] & 6'h3b == _GEN_3921 ? buffer_0_59 : _GEN_1089; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1091 = 2'h0 == read_ptr[1:0] & 6'h3c == _GEN_3921 ? buffer_0_60 : _GEN_1090; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1092 = 2'h0 == read_ptr[1:0] & 6'h3d == _GEN_3921 ? buffer_0_61 : _GEN_1091; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1093 = 2'h0 == read_ptr[1:0] & 6'h3e == _GEN_3921 ? buffer_0_62 : _GEN_1092; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1094 = 2'h0 == read_ptr[1:0] & 6'h3f == _GEN_3921 ? buffer_0_63 : _GEN_1093; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1095 = 2'h1 == read_ptr[1:0] & 5'h0 == _io_out_activate_2_T_4 ? buffer_1_0 : _GEN_1094; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1096 = 2'h1 == read_ptr[1:0] & 5'h1 == _io_out_activate_2_T_4 ? buffer_1_1 : _GEN_1095; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1097 = 2'h1 == read_ptr[1:0] & 5'h2 == _io_out_activate_2_T_4 ? buffer_1_2 : _GEN_1096; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1098 = 2'h1 == read_ptr[1:0] & 5'h3 == _io_out_activate_2_T_4 ? buffer_1_3 : _GEN_1097; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1099 = 2'h1 == read_ptr[1:0] & 5'h4 == _io_out_activate_2_T_4 ? buffer_1_4 : _GEN_1098; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1100 = 2'h1 == read_ptr[1:0] & 5'h5 == _io_out_activate_2_T_4 ? buffer_1_5 : _GEN_1099; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1101 = 2'h1 == read_ptr[1:0] & 5'h6 == _io_out_activate_2_T_4 ? buffer_1_6 : _GEN_1100; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1102 = 2'h1 == read_ptr[1:0] & 5'h7 == _io_out_activate_2_T_4 ? buffer_1_7 : _GEN_1101; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1103 = 2'h1 == read_ptr[1:0] & 5'h8 == _io_out_activate_2_T_4 ? buffer_1_8 : _GEN_1102; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1104 = 2'h1 == read_ptr[1:0] & 5'h9 == _io_out_activate_2_T_4 ? buffer_1_9 : _GEN_1103; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1105 = 2'h1 == read_ptr[1:0] & 5'ha == _io_out_activate_2_T_4 ? buffer_1_10 : _GEN_1104; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1106 = 2'h1 == read_ptr[1:0] & 5'hb == _io_out_activate_2_T_4 ? buffer_1_11 : _GEN_1105; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1107 = 2'h1 == read_ptr[1:0] & 5'hc == _io_out_activate_2_T_4 ? buffer_1_12 : _GEN_1106; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1108 = 2'h1 == read_ptr[1:0] & 5'hd == _io_out_activate_2_T_4 ? buffer_1_13 : _GEN_1107; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1109 = 2'h1 == read_ptr[1:0] & 5'he == _io_out_activate_2_T_4 ? buffer_1_14 : _GEN_1108; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1110 = 2'h1 == read_ptr[1:0] & 5'hf == _io_out_activate_2_T_4 ? buffer_1_15 : _GEN_1109; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1111 = 2'h1 == read_ptr[1:0] & 5'h10 == _io_out_activate_2_T_4 ? buffer_1_16 : _GEN_1110; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1112 = 2'h1 == read_ptr[1:0] & 5'h11 == _io_out_activate_2_T_4 ? buffer_1_17 : _GEN_1111; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1113 = 2'h1 == read_ptr[1:0] & 5'h12 == _io_out_activate_2_T_4 ? buffer_1_18 : _GEN_1112; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1114 = 2'h1 == read_ptr[1:0] & 5'h13 == _io_out_activate_2_T_4 ? buffer_1_19 : _GEN_1113; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1115 = 2'h1 == read_ptr[1:0] & 5'h14 == _io_out_activate_2_T_4 ? buffer_1_20 : _GEN_1114; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1116 = 2'h1 == read_ptr[1:0] & 5'h15 == _io_out_activate_2_T_4 ? buffer_1_21 : _GEN_1115; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1117 = 2'h1 == read_ptr[1:0] & 5'h16 == _io_out_activate_2_T_4 ? buffer_1_22 : _GEN_1116; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1118 = 2'h1 == read_ptr[1:0] & 5'h17 == _io_out_activate_2_T_4 ? buffer_1_23 : _GEN_1117; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1119 = 2'h1 == read_ptr[1:0] & 5'h18 == _io_out_activate_2_T_4 ? buffer_1_24 : _GEN_1118; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1120 = 2'h1 == read_ptr[1:0] & 5'h19 == _io_out_activate_2_T_4 ? buffer_1_25 : _GEN_1119; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1121 = 2'h1 == read_ptr[1:0] & 5'h1a == _io_out_activate_2_T_4 ? buffer_1_26 : _GEN_1120; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1122 = 2'h1 == read_ptr[1:0] & 5'h1b == _io_out_activate_2_T_4 ? buffer_1_27 : _GEN_1121; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1123 = 2'h1 == read_ptr[1:0] & 5'h1c == _io_out_activate_2_T_4 ? buffer_1_28 : _GEN_1122; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1124 = 2'h1 == read_ptr[1:0] & 5'h1d == _io_out_activate_2_T_4 ? buffer_1_29 : _GEN_1123; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1125 = 2'h1 == read_ptr[1:0] & 5'h1e == _io_out_activate_2_T_4 ? buffer_1_30 : _GEN_1124; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1126 = 2'h1 == read_ptr[1:0] & 5'h1f == _io_out_activate_2_T_4 ? buffer_1_31 : _GEN_1125; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1127 = 2'h1 == read_ptr[1:0] & 6'h20 == _GEN_3921 ? buffer_1_32 : _GEN_1126; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1128 = 2'h1 == read_ptr[1:0] & 6'h21 == _GEN_3921 ? buffer_1_33 : _GEN_1127; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1129 = 2'h1 == read_ptr[1:0] & 6'h22 == _GEN_3921 ? buffer_1_34 : _GEN_1128; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1130 = 2'h1 == read_ptr[1:0] & 6'h23 == _GEN_3921 ? buffer_1_35 : _GEN_1129; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1131 = 2'h1 == read_ptr[1:0] & 6'h24 == _GEN_3921 ? buffer_1_36 : _GEN_1130; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1132 = 2'h1 == read_ptr[1:0] & 6'h25 == _GEN_3921 ? buffer_1_37 : _GEN_1131; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1133 = 2'h1 == read_ptr[1:0] & 6'h26 == _GEN_3921 ? buffer_1_38 : _GEN_1132; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1134 = 2'h1 == read_ptr[1:0] & 6'h27 == _GEN_3921 ? buffer_1_39 : _GEN_1133; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1135 = 2'h1 == read_ptr[1:0] & 6'h28 == _GEN_3921 ? buffer_1_40 : _GEN_1134; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1136 = 2'h1 == read_ptr[1:0] & 6'h29 == _GEN_3921 ? buffer_1_41 : _GEN_1135; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1137 = 2'h1 == read_ptr[1:0] & 6'h2a == _GEN_3921 ? buffer_1_42 : _GEN_1136; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1138 = 2'h1 == read_ptr[1:0] & 6'h2b == _GEN_3921 ? buffer_1_43 : _GEN_1137; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1139 = 2'h1 == read_ptr[1:0] & 6'h2c == _GEN_3921 ? buffer_1_44 : _GEN_1138; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1140 = 2'h1 == read_ptr[1:0] & 6'h2d == _GEN_3921 ? buffer_1_45 : _GEN_1139; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1141 = 2'h1 == read_ptr[1:0] & 6'h2e == _GEN_3921 ? buffer_1_46 : _GEN_1140; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1142 = 2'h1 == read_ptr[1:0] & 6'h2f == _GEN_3921 ? buffer_1_47 : _GEN_1141; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1143 = 2'h1 == read_ptr[1:0] & 6'h30 == _GEN_3921 ? buffer_1_48 : _GEN_1142; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1144 = 2'h1 == read_ptr[1:0] & 6'h31 == _GEN_3921 ? buffer_1_49 : _GEN_1143; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1145 = 2'h1 == read_ptr[1:0] & 6'h32 == _GEN_3921 ? buffer_1_50 : _GEN_1144; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1146 = 2'h1 == read_ptr[1:0] & 6'h33 == _GEN_3921 ? buffer_1_51 : _GEN_1145; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1147 = 2'h1 == read_ptr[1:0] & 6'h34 == _GEN_3921 ? buffer_1_52 : _GEN_1146; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1148 = 2'h1 == read_ptr[1:0] & 6'h35 == _GEN_3921 ? buffer_1_53 : _GEN_1147; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1149 = 2'h1 == read_ptr[1:0] & 6'h36 == _GEN_3921 ? buffer_1_54 : _GEN_1148; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1150 = 2'h1 == read_ptr[1:0] & 6'h37 == _GEN_3921 ? buffer_1_55 : _GEN_1149; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1151 = 2'h1 == read_ptr[1:0] & 6'h38 == _GEN_3921 ? buffer_1_56 : _GEN_1150; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1152 = 2'h1 == read_ptr[1:0] & 6'h39 == _GEN_3921 ? buffer_1_57 : _GEN_1151; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1153 = 2'h1 == read_ptr[1:0] & 6'h3a == _GEN_3921 ? buffer_1_58 : _GEN_1152; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1154 = 2'h1 == read_ptr[1:0] & 6'h3b == _GEN_3921 ? buffer_1_59 : _GEN_1153; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1155 = 2'h1 == read_ptr[1:0] & 6'h3c == _GEN_3921 ? buffer_1_60 : _GEN_1154; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1156 = 2'h1 == read_ptr[1:0] & 6'h3d == _GEN_3921 ? buffer_1_61 : _GEN_1155; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1157 = 2'h1 == read_ptr[1:0] & 6'h3e == _GEN_3921 ? buffer_1_62 : _GEN_1156; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1158 = 2'h1 == read_ptr[1:0] & 6'h3f == _GEN_3921 ? buffer_1_63 : _GEN_1157; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1159 = 2'h2 == read_ptr[1:0] & 5'h0 == _io_out_activate_2_T_4 ? buffer_2_0 : _GEN_1158; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1160 = 2'h2 == read_ptr[1:0] & 5'h1 == _io_out_activate_2_T_4 ? buffer_2_1 : _GEN_1159; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1161 = 2'h2 == read_ptr[1:0] & 5'h2 == _io_out_activate_2_T_4 ? buffer_2_2 : _GEN_1160; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1162 = 2'h2 == read_ptr[1:0] & 5'h3 == _io_out_activate_2_T_4 ? buffer_2_3 : _GEN_1161; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1163 = 2'h2 == read_ptr[1:0] & 5'h4 == _io_out_activate_2_T_4 ? buffer_2_4 : _GEN_1162; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1164 = 2'h2 == read_ptr[1:0] & 5'h5 == _io_out_activate_2_T_4 ? buffer_2_5 : _GEN_1163; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1165 = 2'h2 == read_ptr[1:0] & 5'h6 == _io_out_activate_2_T_4 ? buffer_2_6 : _GEN_1164; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1166 = 2'h2 == read_ptr[1:0] & 5'h7 == _io_out_activate_2_T_4 ? buffer_2_7 : _GEN_1165; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1167 = 2'h2 == read_ptr[1:0] & 5'h8 == _io_out_activate_2_T_4 ? buffer_2_8 : _GEN_1166; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1168 = 2'h2 == read_ptr[1:0] & 5'h9 == _io_out_activate_2_T_4 ? buffer_2_9 : _GEN_1167; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1169 = 2'h2 == read_ptr[1:0] & 5'ha == _io_out_activate_2_T_4 ? buffer_2_10 : _GEN_1168; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1170 = 2'h2 == read_ptr[1:0] & 5'hb == _io_out_activate_2_T_4 ? buffer_2_11 : _GEN_1169; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1171 = 2'h2 == read_ptr[1:0] & 5'hc == _io_out_activate_2_T_4 ? buffer_2_12 : _GEN_1170; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1172 = 2'h2 == read_ptr[1:0] & 5'hd == _io_out_activate_2_T_4 ? buffer_2_13 : _GEN_1171; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1173 = 2'h2 == read_ptr[1:0] & 5'he == _io_out_activate_2_T_4 ? buffer_2_14 : _GEN_1172; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1174 = 2'h2 == read_ptr[1:0] & 5'hf == _io_out_activate_2_T_4 ? buffer_2_15 : _GEN_1173; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1175 = 2'h2 == read_ptr[1:0] & 5'h10 == _io_out_activate_2_T_4 ? buffer_2_16 : _GEN_1174; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1176 = 2'h2 == read_ptr[1:0] & 5'h11 == _io_out_activate_2_T_4 ? buffer_2_17 : _GEN_1175; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1177 = 2'h2 == read_ptr[1:0] & 5'h12 == _io_out_activate_2_T_4 ? buffer_2_18 : _GEN_1176; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1178 = 2'h2 == read_ptr[1:0] & 5'h13 == _io_out_activate_2_T_4 ? buffer_2_19 : _GEN_1177; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1179 = 2'h2 == read_ptr[1:0] & 5'h14 == _io_out_activate_2_T_4 ? buffer_2_20 : _GEN_1178; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1180 = 2'h2 == read_ptr[1:0] & 5'h15 == _io_out_activate_2_T_4 ? buffer_2_21 : _GEN_1179; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1181 = 2'h2 == read_ptr[1:0] & 5'h16 == _io_out_activate_2_T_4 ? buffer_2_22 : _GEN_1180; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1182 = 2'h2 == read_ptr[1:0] & 5'h17 == _io_out_activate_2_T_4 ? buffer_2_23 : _GEN_1181; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1183 = 2'h2 == read_ptr[1:0] & 5'h18 == _io_out_activate_2_T_4 ? buffer_2_24 : _GEN_1182; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1184 = 2'h2 == read_ptr[1:0] & 5'h19 == _io_out_activate_2_T_4 ? buffer_2_25 : _GEN_1183; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1185 = 2'h2 == read_ptr[1:0] & 5'h1a == _io_out_activate_2_T_4 ? buffer_2_26 : _GEN_1184; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1186 = 2'h2 == read_ptr[1:0] & 5'h1b == _io_out_activate_2_T_4 ? buffer_2_27 : _GEN_1185; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1187 = 2'h2 == read_ptr[1:0] & 5'h1c == _io_out_activate_2_T_4 ? buffer_2_28 : _GEN_1186; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1188 = 2'h2 == read_ptr[1:0] & 5'h1d == _io_out_activate_2_T_4 ? buffer_2_29 : _GEN_1187; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1189 = 2'h2 == read_ptr[1:0] & 5'h1e == _io_out_activate_2_T_4 ? buffer_2_30 : _GEN_1188; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1190 = 2'h2 == read_ptr[1:0] & 5'h1f == _io_out_activate_2_T_4 ? buffer_2_31 : _GEN_1189; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1191 = 2'h2 == read_ptr[1:0] & 6'h20 == _GEN_3921 ? buffer_2_32 : _GEN_1190; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1192 = 2'h2 == read_ptr[1:0] & 6'h21 == _GEN_3921 ? buffer_2_33 : _GEN_1191; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1193 = 2'h2 == read_ptr[1:0] & 6'h22 == _GEN_3921 ? buffer_2_34 : _GEN_1192; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1194 = 2'h2 == read_ptr[1:0] & 6'h23 == _GEN_3921 ? buffer_2_35 : _GEN_1193; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1195 = 2'h2 == read_ptr[1:0] & 6'h24 == _GEN_3921 ? buffer_2_36 : _GEN_1194; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1196 = 2'h2 == read_ptr[1:0] & 6'h25 == _GEN_3921 ? buffer_2_37 : _GEN_1195; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1197 = 2'h2 == read_ptr[1:0] & 6'h26 == _GEN_3921 ? buffer_2_38 : _GEN_1196; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1198 = 2'h2 == read_ptr[1:0] & 6'h27 == _GEN_3921 ? buffer_2_39 : _GEN_1197; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1199 = 2'h2 == read_ptr[1:0] & 6'h28 == _GEN_3921 ? buffer_2_40 : _GEN_1198; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1200 = 2'h2 == read_ptr[1:0] & 6'h29 == _GEN_3921 ? buffer_2_41 : _GEN_1199; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1201 = 2'h2 == read_ptr[1:0] & 6'h2a == _GEN_3921 ? buffer_2_42 : _GEN_1200; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1202 = 2'h2 == read_ptr[1:0] & 6'h2b == _GEN_3921 ? buffer_2_43 : _GEN_1201; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1203 = 2'h2 == read_ptr[1:0] & 6'h2c == _GEN_3921 ? buffer_2_44 : _GEN_1202; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1204 = 2'h2 == read_ptr[1:0] & 6'h2d == _GEN_3921 ? buffer_2_45 : _GEN_1203; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1205 = 2'h2 == read_ptr[1:0] & 6'h2e == _GEN_3921 ? buffer_2_46 : _GEN_1204; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1206 = 2'h2 == read_ptr[1:0] & 6'h2f == _GEN_3921 ? buffer_2_47 : _GEN_1205; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1207 = 2'h2 == read_ptr[1:0] & 6'h30 == _GEN_3921 ? buffer_2_48 : _GEN_1206; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1208 = 2'h2 == read_ptr[1:0] & 6'h31 == _GEN_3921 ? buffer_2_49 : _GEN_1207; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1209 = 2'h2 == read_ptr[1:0] & 6'h32 == _GEN_3921 ? buffer_2_50 : _GEN_1208; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1210 = 2'h2 == read_ptr[1:0] & 6'h33 == _GEN_3921 ? buffer_2_51 : _GEN_1209; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1211 = 2'h2 == read_ptr[1:0] & 6'h34 == _GEN_3921 ? buffer_2_52 : _GEN_1210; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1212 = 2'h2 == read_ptr[1:0] & 6'h35 == _GEN_3921 ? buffer_2_53 : _GEN_1211; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1213 = 2'h2 == read_ptr[1:0] & 6'h36 == _GEN_3921 ? buffer_2_54 : _GEN_1212; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1214 = 2'h2 == read_ptr[1:0] & 6'h37 == _GEN_3921 ? buffer_2_55 : _GEN_1213; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1215 = 2'h2 == read_ptr[1:0] & 6'h38 == _GEN_3921 ? buffer_2_56 : _GEN_1214; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1216 = 2'h2 == read_ptr[1:0] & 6'h39 == _GEN_3921 ? buffer_2_57 : _GEN_1215; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1217 = 2'h2 == read_ptr[1:0] & 6'h3a == _GEN_3921 ? buffer_2_58 : _GEN_1216; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1218 = 2'h2 == read_ptr[1:0] & 6'h3b == _GEN_3921 ? buffer_2_59 : _GEN_1217; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1219 = 2'h2 == read_ptr[1:0] & 6'h3c == _GEN_3921 ? buffer_2_60 : _GEN_1218; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1220 = 2'h2 == read_ptr[1:0] & 6'h3d == _GEN_3921 ? buffer_2_61 : _GEN_1219; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1221 = 2'h2 == read_ptr[1:0] & 6'h3e == _GEN_3921 ? buffer_2_62 : _GEN_1220; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1222 = 2'h2 == read_ptr[1:0] & 6'h3f == _GEN_3921 ? buffer_2_63 : _GEN_1221; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1223 = 2'h3 == read_ptr[1:0] & 5'h0 == _io_out_activate_2_T_4 ? buffer_3_0 : _GEN_1222; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1224 = 2'h3 == read_ptr[1:0] & 5'h1 == _io_out_activate_2_T_4 ? buffer_3_1 : _GEN_1223; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1225 = 2'h3 == read_ptr[1:0] & 5'h2 == _io_out_activate_2_T_4 ? buffer_3_2 : _GEN_1224; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1226 = 2'h3 == read_ptr[1:0] & 5'h3 == _io_out_activate_2_T_4 ? buffer_3_3 : _GEN_1225; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1227 = 2'h3 == read_ptr[1:0] & 5'h4 == _io_out_activate_2_T_4 ? buffer_3_4 : _GEN_1226; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1228 = 2'h3 == read_ptr[1:0] & 5'h5 == _io_out_activate_2_T_4 ? buffer_3_5 : _GEN_1227; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1229 = 2'h3 == read_ptr[1:0] & 5'h6 == _io_out_activate_2_T_4 ? buffer_3_6 : _GEN_1228; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1230 = 2'h3 == read_ptr[1:0] & 5'h7 == _io_out_activate_2_T_4 ? buffer_3_7 : _GEN_1229; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1231 = 2'h3 == read_ptr[1:0] & 5'h8 == _io_out_activate_2_T_4 ? buffer_3_8 : _GEN_1230; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1232 = 2'h3 == read_ptr[1:0] & 5'h9 == _io_out_activate_2_T_4 ? buffer_3_9 : _GEN_1231; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1233 = 2'h3 == read_ptr[1:0] & 5'ha == _io_out_activate_2_T_4 ? buffer_3_10 : _GEN_1232; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1234 = 2'h3 == read_ptr[1:0] & 5'hb == _io_out_activate_2_T_4 ? buffer_3_11 : _GEN_1233; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1235 = 2'h3 == read_ptr[1:0] & 5'hc == _io_out_activate_2_T_4 ? buffer_3_12 : _GEN_1234; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1236 = 2'h3 == read_ptr[1:0] & 5'hd == _io_out_activate_2_T_4 ? buffer_3_13 : _GEN_1235; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1237 = 2'h3 == read_ptr[1:0] & 5'he == _io_out_activate_2_T_4 ? buffer_3_14 : _GEN_1236; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1238 = 2'h3 == read_ptr[1:0] & 5'hf == _io_out_activate_2_T_4 ? buffer_3_15 : _GEN_1237; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1239 = 2'h3 == read_ptr[1:0] & 5'h10 == _io_out_activate_2_T_4 ? buffer_3_16 : _GEN_1238; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1240 = 2'h3 == read_ptr[1:0] & 5'h11 == _io_out_activate_2_T_4 ? buffer_3_17 : _GEN_1239; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1241 = 2'h3 == read_ptr[1:0] & 5'h12 == _io_out_activate_2_T_4 ? buffer_3_18 : _GEN_1240; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1242 = 2'h3 == read_ptr[1:0] & 5'h13 == _io_out_activate_2_T_4 ? buffer_3_19 : _GEN_1241; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1243 = 2'h3 == read_ptr[1:0] & 5'h14 == _io_out_activate_2_T_4 ? buffer_3_20 : _GEN_1242; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1244 = 2'h3 == read_ptr[1:0] & 5'h15 == _io_out_activate_2_T_4 ? buffer_3_21 : _GEN_1243; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1245 = 2'h3 == read_ptr[1:0] & 5'h16 == _io_out_activate_2_T_4 ? buffer_3_22 : _GEN_1244; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1246 = 2'h3 == read_ptr[1:0] & 5'h17 == _io_out_activate_2_T_4 ? buffer_3_23 : _GEN_1245; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1247 = 2'h3 == read_ptr[1:0] & 5'h18 == _io_out_activate_2_T_4 ? buffer_3_24 : _GEN_1246; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1248 = 2'h3 == read_ptr[1:0] & 5'h19 == _io_out_activate_2_T_4 ? buffer_3_25 : _GEN_1247; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1249 = 2'h3 == read_ptr[1:0] & 5'h1a == _io_out_activate_2_T_4 ? buffer_3_26 : _GEN_1248; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1250 = 2'h3 == read_ptr[1:0] & 5'h1b == _io_out_activate_2_T_4 ? buffer_3_27 : _GEN_1249; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1251 = 2'h3 == read_ptr[1:0] & 5'h1c == _io_out_activate_2_T_4 ? buffer_3_28 : _GEN_1250; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1252 = 2'h3 == read_ptr[1:0] & 5'h1d == _io_out_activate_2_T_4 ? buffer_3_29 : _GEN_1251; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1253 = 2'h3 == read_ptr[1:0] & 5'h1e == _io_out_activate_2_T_4 ? buffer_3_30 : _GEN_1252; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1254 = 2'h3 == read_ptr[1:0] & 5'h1f == _io_out_activate_2_T_4 ? buffer_3_31 : _GEN_1253; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1255 = 2'h3 == read_ptr[1:0] & 6'h20 == _GEN_3921 ? buffer_3_32 : _GEN_1254; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1256 = 2'h3 == read_ptr[1:0] & 6'h21 == _GEN_3921 ? buffer_3_33 : _GEN_1255; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1257 = 2'h3 == read_ptr[1:0] & 6'h22 == _GEN_3921 ? buffer_3_34 : _GEN_1256; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1258 = 2'h3 == read_ptr[1:0] & 6'h23 == _GEN_3921 ? buffer_3_35 : _GEN_1257; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1259 = 2'h3 == read_ptr[1:0] & 6'h24 == _GEN_3921 ? buffer_3_36 : _GEN_1258; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1260 = 2'h3 == read_ptr[1:0] & 6'h25 == _GEN_3921 ? buffer_3_37 : _GEN_1259; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1261 = 2'h3 == read_ptr[1:0] & 6'h26 == _GEN_3921 ? buffer_3_38 : _GEN_1260; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1262 = 2'h3 == read_ptr[1:0] & 6'h27 == _GEN_3921 ? buffer_3_39 : _GEN_1261; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1263 = 2'h3 == read_ptr[1:0] & 6'h28 == _GEN_3921 ? buffer_3_40 : _GEN_1262; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1264 = 2'h3 == read_ptr[1:0] & 6'h29 == _GEN_3921 ? buffer_3_41 : _GEN_1263; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1265 = 2'h3 == read_ptr[1:0] & 6'h2a == _GEN_3921 ? buffer_3_42 : _GEN_1264; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1266 = 2'h3 == read_ptr[1:0] & 6'h2b == _GEN_3921 ? buffer_3_43 : _GEN_1265; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1267 = 2'h3 == read_ptr[1:0] & 6'h2c == _GEN_3921 ? buffer_3_44 : _GEN_1266; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1268 = 2'h3 == read_ptr[1:0] & 6'h2d == _GEN_3921 ? buffer_3_45 : _GEN_1267; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1269 = 2'h3 == read_ptr[1:0] & 6'h2e == _GEN_3921 ? buffer_3_46 : _GEN_1268; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1270 = 2'h3 == read_ptr[1:0] & 6'h2f == _GEN_3921 ? buffer_3_47 : _GEN_1269; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1271 = 2'h3 == read_ptr[1:0] & 6'h30 == _GEN_3921 ? buffer_3_48 : _GEN_1270; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1272 = 2'h3 == read_ptr[1:0] & 6'h31 == _GEN_3921 ? buffer_3_49 : _GEN_1271; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1273 = 2'h3 == read_ptr[1:0] & 6'h32 == _GEN_3921 ? buffer_3_50 : _GEN_1272; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1274 = 2'h3 == read_ptr[1:0] & 6'h33 == _GEN_3921 ? buffer_3_51 : _GEN_1273; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1275 = 2'h3 == read_ptr[1:0] & 6'h34 == _GEN_3921 ? buffer_3_52 : _GEN_1274; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1276 = 2'h3 == read_ptr[1:0] & 6'h35 == _GEN_3921 ? buffer_3_53 : _GEN_1275; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1277 = 2'h3 == read_ptr[1:0] & 6'h36 == _GEN_3921 ? buffer_3_54 : _GEN_1276; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1278 = 2'h3 == read_ptr[1:0] & 6'h37 == _GEN_3921 ? buffer_3_55 : _GEN_1277; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1279 = 2'h3 == read_ptr[1:0] & 6'h38 == _GEN_3921 ? buffer_3_56 : _GEN_1278; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1280 = 2'h3 == read_ptr[1:0] & 6'h39 == _GEN_3921 ? buffer_3_57 : _GEN_1279; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1281 = 2'h3 == read_ptr[1:0] & 6'h3a == _GEN_3921 ? buffer_3_58 : _GEN_1280; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1282 = 2'h3 == read_ptr[1:0] & 6'h3b == _GEN_3921 ? buffer_3_59 : _GEN_1281; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1283 = 2'h3 == read_ptr[1:0] & 6'h3c == _GEN_3921 ? buffer_3_60 : _GEN_1282; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1284 = 2'h3 == read_ptr[1:0] & 6'h3d == _GEN_3921 ? buffer_3_61 : _GEN_1283; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1285 = 2'h3 == read_ptr[1:0] & 6'h3e == _GEN_3921 ? buffer_3_62 : _GEN_1284; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1286 = 2'h3 == read_ptr[1:0] & 6'h3f == _GEN_3921 ? buffer_3_63 : _GEN_1285; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1287 = 5'h2 < flow_ptr & flow_ptr <= 5'ha ? _GEN_1286 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [4:0] _io_out_activate_3_T_2 = 5'h18 + flow_ptr; // @[Activation_Buffer.scala 76:88]
  wire [4:0] _io_out_activate_3_T_4 = _io_out_activate_3_T_2 - 5'h4; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_1289 = 2'h0 == read_ptr[1:0] & 5'h1 == _io_out_activate_3_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1290 = 2'h0 == read_ptr[1:0] & 5'h2 == _io_out_activate_3_T_4 ? buffer_0_2 : _GEN_1289; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1291 = 2'h0 == read_ptr[1:0] & 5'h3 == _io_out_activate_3_T_4 ? buffer_0_3 : _GEN_1290; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1292 = 2'h0 == read_ptr[1:0] & 5'h4 == _io_out_activate_3_T_4 ? buffer_0_4 : _GEN_1291; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1293 = 2'h0 == read_ptr[1:0] & 5'h5 == _io_out_activate_3_T_4 ? buffer_0_5 : _GEN_1292; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1294 = 2'h0 == read_ptr[1:0] & 5'h6 == _io_out_activate_3_T_4 ? buffer_0_6 : _GEN_1293; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1295 = 2'h0 == read_ptr[1:0] & 5'h7 == _io_out_activate_3_T_4 ? buffer_0_7 : _GEN_1294; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1296 = 2'h0 == read_ptr[1:0] & 5'h8 == _io_out_activate_3_T_4 ? buffer_0_8 : _GEN_1295; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1297 = 2'h0 == read_ptr[1:0] & 5'h9 == _io_out_activate_3_T_4 ? buffer_0_9 : _GEN_1296; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1298 = 2'h0 == read_ptr[1:0] & 5'ha == _io_out_activate_3_T_4 ? buffer_0_10 : _GEN_1297; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1299 = 2'h0 == read_ptr[1:0] & 5'hb == _io_out_activate_3_T_4 ? buffer_0_11 : _GEN_1298; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1300 = 2'h0 == read_ptr[1:0] & 5'hc == _io_out_activate_3_T_4 ? buffer_0_12 : _GEN_1299; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1301 = 2'h0 == read_ptr[1:0] & 5'hd == _io_out_activate_3_T_4 ? buffer_0_13 : _GEN_1300; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1302 = 2'h0 == read_ptr[1:0] & 5'he == _io_out_activate_3_T_4 ? buffer_0_14 : _GEN_1301; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1303 = 2'h0 == read_ptr[1:0] & 5'hf == _io_out_activate_3_T_4 ? buffer_0_15 : _GEN_1302; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1304 = 2'h0 == read_ptr[1:0] & 5'h10 == _io_out_activate_3_T_4 ? buffer_0_16 : _GEN_1303; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1305 = 2'h0 == read_ptr[1:0] & 5'h11 == _io_out_activate_3_T_4 ? buffer_0_17 : _GEN_1304; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1306 = 2'h0 == read_ptr[1:0] & 5'h12 == _io_out_activate_3_T_4 ? buffer_0_18 : _GEN_1305; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1307 = 2'h0 == read_ptr[1:0] & 5'h13 == _io_out_activate_3_T_4 ? buffer_0_19 : _GEN_1306; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1308 = 2'h0 == read_ptr[1:0] & 5'h14 == _io_out_activate_3_T_4 ? buffer_0_20 : _GEN_1307; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1309 = 2'h0 == read_ptr[1:0] & 5'h15 == _io_out_activate_3_T_4 ? buffer_0_21 : _GEN_1308; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1310 = 2'h0 == read_ptr[1:0] & 5'h16 == _io_out_activate_3_T_4 ? buffer_0_22 : _GEN_1309; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1311 = 2'h0 == read_ptr[1:0] & 5'h17 == _io_out_activate_3_T_4 ? buffer_0_23 : _GEN_1310; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1312 = 2'h0 == read_ptr[1:0] & 5'h18 == _io_out_activate_3_T_4 ? buffer_0_24 : _GEN_1311; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1313 = 2'h0 == read_ptr[1:0] & 5'h19 == _io_out_activate_3_T_4 ? buffer_0_25 : _GEN_1312; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1314 = 2'h0 == read_ptr[1:0] & 5'h1a == _io_out_activate_3_T_4 ? buffer_0_26 : _GEN_1313; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1315 = 2'h0 == read_ptr[1:0] & 5'h1b == _io_out_activate_3_T_4 ? buffer_0_27 : _GEN_1314; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1316 = 2'h0 == read_ptr[1:0] & 5'h1c == _io_out_activate_3_T_4 ? buffer_0_28 : _GEN_1315; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1317 = 2'h0 == read_ptr[1:0] & 5'h1d == _io_out_activate_3_T_4 ? buffer_0_29 : _GEN_1316; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1318 = 2'h0 == read_ptr[1:0] & 5'h1e == _io_out_activate_3_T_4 ? buffer_0_30 : _GEN_1317; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1319 = 2'h0 == read_ptr[1:0] & 5'h1f == _io_out_activate_3_T_4 ? buffer_0_31 : _GEN_1318; // @[Activation_Buffer.scala 76:{28,28}]
  wire [5:0] _GEN_4559 = {{1'd0}, _io_out_activate_3_T_4}; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1320 = 2'h0 == read_ptr[1:0] & 6'h20 == _GEN_4559 ? buffer_0_32 : _GEN_1319; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1321 = 2'h0 == read_ptr[1:0] & 6'h21 == _GEN_4559 ? buffer_0_33 : _GEN_1320; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1322 = 2'h0 == read_ptr[1:0] & 6'h22 == _GEN_4559 ? buffer_0_34 : _GEN_1321; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1323 = 2'h0 == read_ptr[1:0] & 6'h23 == _GEN_4559 ? buffer_0_35 : _GEN_1322; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1324 = 2'h0 == read_ptr[1:0] & 6'h24 == _GEN_4559 ? buffer_0_36 : _GEN_1323; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1325 = 2'h0 == read_ptr[1:0] & 6'h25 == _GEN_4559 ? buffer_0_37 : _GEN_1324; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1326 = 2'h0 == read_ptr[1:0] & 6'h26 == _GEN_4559 ? buffer_0_38 : _GEN_1325; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1327 = 2'h0 == read_ptr[1:0] & 6'h27 == _GEN_4559 ? buffer_0_39 : _GEN_1326; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1328 = 2'h0 == read_ptr[1:0] & 6'h28 == _GEN_4559 ? buffer_0_40 : _GEN_1327; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1329 = 2'h0 == read_ptr[1:0] & 6'h29 == _GEN_4559 ? buffer_0_41 : _GEN_1328; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1330 = 2'h0 == read_ptr[1:0] & 6'h2a == _GEN_4559 ? buffer_0_42 : _GEN_1329; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1331 = 2'h0 == read_ptr[1:0] & 6'h2b == _GEN_4559 ? buffer_0_43 : _GEN_1330; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1332 = 2'h0 == read_ptr[1:0] & 6'h2c == _GEN_4559 ? buffer_0_44 : _GEN_1331; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1333 = 2'h0 == read_ptr[1:0] & 6'h2d == _GEN_4559 ? buffer_0_45 : _GEN_1332; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1334 = 2'h0 == read_ptr[1:0] & 6'h2e == _GEN_4559 ? buffer_0_46 : _GEN_1333; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1335 = 2'h0 == read_ptr[1:0] & 6'h2f == _GEN_4559 ? buffer_0_47 : _GEN_1334; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1336 = 2'h0 == read_ptr[1:0] & 6'h30 == _GEN_4559 ? buffer_0_48 : _GEN_1335; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1337 = 2'h0 == read_ptr[1:0] & 6'h31 == _GEN_4559 ? buffer_0_49 : _GEN_1336; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1338 = 2'h0 == read_ptr[1:0] & 6'h32 == _GEN_4559 ? buffer_0_50 : _GEN_1337; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1339 = 2'h0 == read_ptr[1:0] & 6'h33 == _GEN_4559 ? buffer_0_51 : _GEN_1338; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1340 = 2'h0 == read_ptr[1:0] & 6'h34 == _GEN_4559 ? buffer_0_52 : _GEN_1339; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1341 = 2'h0 == read_ptr[1:0] & 6'h35 == _GEN_4559 ? buffer_0_53 : _GEN_1340; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1342 = 2'h0 == read_ptr[1:0] & 6'h36 == _GEN_4559 ? buffer_0_54 : _GEN_1341; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1343 = 2'h0 == read_ptr[1:0] & 6'h37 == _GEN_4559 ? buffer_0_55 : _GEN_1342; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1344 = 2'h0 == read_ptr[1:0] & 6'h38 == _GEN_4559 ? buffer_0_56 : _GEN_1343; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1345 = 2'h0 == read_ptr[1:0] & 6'h39 == _GEN_4559 ? buffer_0_57 : _GEN_1344; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1346 = 2'h0 == read_ptr[1:0] & 6'h3a == _GEN_4559 ? buffer_0_58 : _GEN_1345; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1347 = 2'h0 == read_ptr[1:0] & 6'h3b == _GEN_4559 ? buffer_0_59 : _GEN_1346; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1348 = 2'h0 == read_ptr[1:0] & 6'h3c == _GEN_4559 ? buffer_0_60 : _GEN_1347; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1349 = 2'h0 == read_ptr[1:0] & 6'h3d == _GEN_4559 ? buffer_0_61 : _GEN_1348; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1350 = 2'h0 == read_ptr[1:0] & 6'h3e == _GEN_4559 ? buffer_0_62 : _GEN_1349; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1351 = 2'h0 == read_ptr[1:0] & 6'h3f == _GEN_4559 ? buffer_0_63 : _GEN_1350; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1352 = 2'h1 == read_ptr[1:0] & 5'h0 == _io_out_activate_3_T_4 ? buffer_1_0 : _GEN_1351; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1353 = 2'h1 == read_ptr[1:0] & 5'h1 == _io_out_activate_3_T_4 ? buffer_1_1 : _GEN_1352; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1354 = 2'h1 == read_ptr[1:0] & 5'h2 == _io_out_activate_3_T_4 ? buffer_1_2 : _GEN_1353; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1355 = 2'h1 == read_ptr[1:0] & 5'h3 == _io_out_activate_3_T_4 ? buffer_1_3 : _GEN_1354; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1356 = 2'h1 == read_ptr[1:0] & 5'h4 == _io_out_activate_3_T_4 ? buffer_1_4 : _GEN_1355; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1357 = 2'h1 == read_ptr[1:0] & 5'h5 == _io_out_activate_3_T_4 ? buffer_1_5 : _GEN_1356; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1358 = 2'h1 == read_ptr[1:0] & 5'h6 == _io_out_activate_3_T_4 ? buffer_1_6 : _GEN_1357; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1359 = 2'h1 == read_ptr[1:0] & 5'h7 == _io_out_activate_3_T_4 ? buffer_1_7 : _GEN_1358; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1360 = 2'h1 == read_ptr[1:0] & 5'h8 == _io_out_activate_3_T_4 ? buffer_1_8 : _GEN_1359; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1361 = 2'h1 == read_ptr[1:0] & 5'h9 == _io_out_activate_3_T_4 ? buffer_1_9 : _GEN_1360; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1362 = 2'h1 == read_ptr[1:0] & 5'ha == _io_out_activate_3_T_4 ? buffer_1_10 : _GEN_1361; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1363 = 2'h1 == read_ptr[1:0] & 5'hb == _io_out_activate_3_T_4 ? buffer_1_11 : _GEN_1362; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1364 = 2'h1 == read_ptr[1:0] & 5'hc == _io_out_activate_3_T_4 ? buffer_1_12 : _GEN_1363; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1365 = 2'h1 == read_ptr[1:0] & 5'hd == _io_out_activate_3_T_4 ? buffer_1_13 : _GEN_1364; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1366 = 2'h1 == read_ptr[1:0] & 5'he == _io_out_activate_3_T_4 ? buffer_1_14 : _GEN_1365; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1367 = 2'h1 == read_ptr[1:0] & 5'hf == _io_out_activate_3_T_4 ? buffer_1_15 : _GEN_1366; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1368 = 2'h1 == read_ptr[1:0] & 5'h10 == _io_out_activate_3_T_4 ? buffer_1_16 : _GEN_1367; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1369 = 2'h1 == read_ptr[1:0] & 5'h11 == _io_out_activate_3_T_4 ? buffer_1_17 : _GEN_1368; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1370 = 2'h1 == read_ptr[1:0] & 5'h12 == _io_out_activate_3_T_4 ? buffer_1_18 : _GEN_1369; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1371 = 2'h1 == read_ptr[1:0] & 5'h13 == _io_out_activate_3_T_4 ? buffer_1_19 : _GEN_1370; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1372 = 2'h1 == read_ptr[1:0] & 5'h14 == _io_out_activate_3_T_4 ? buffer_1_20 : _GEN_1371; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1373 = 2'h1 == read_ptr[1:0] & 5'h15 == _io_out_activate_3_T_4 ? buffer_1_21 : _GEN_1372; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1374 = 2'h1 == read_ptr[1:0] & 5'h16 == _io_out_activate_3_T_4 ? buffer_1_22 : _GEN_1373; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1375 = 2'h1 == read_ptr[1:0] & 5'h17 == _io_out_activate_3_T_4 ? buffer_1_23 : _GEN_1374; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1376 = 2'h1 == read_ptr[1:0] & 5'h18 == _io_out_activate_3_T_4 ? buffer_1_24 : _GEN_1375; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1377 = 2'h1 == read_ptr[1:0] & 5'h19 == _io_out_activate_3_T_4 ? buffer_1_25 : _GEN_1376; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1378 = 2'h1 == read_ptr[1:0] & 5'h1a == _io_out_activate_3_T_4 ? buffer_1_26 : _GEN_1377; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1379 = 2'h1 == read_ptr[1:0] & 5'h1b == _io_out_activate_3_T_4 ? buffer_1_27 : _GEN_1378; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1380 = 2'h1 == read_ptr[1:0] & 5'h1c == _io_out_activate_3_T_4 ? buffer_1_28 : _GEN_1379; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1381 = 2'h1 == read_ptr[1:0] & 5'h1d == _io_out_activate_3_T_4 ? buffer_1_29 : _GEN_1380; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1382 = 2'h1 == read_ptr[1:0] & 5'h1e == _io_out_activate_3_T_4 ? buffer_1_30 : _GEN_1381; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1383 = 2'h1 == read_ptr[1:0] & 5'h1f == _io_out_activate_3_T_4 ? buffer_1_31 : _GEN_1382; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1384 = 2'h1 == read_ptr[1:0] & 6'h20 == _GEN_4559 ? buffer_1_32 : _GEN_1383; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1385 = 2'h1 == read_ptr[1:0] & 6'h21 == _GEN_4559 ? buffer_1_33 : _GEN_1384; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1386 = 2'h1 == read_ptr[1:0] & 6'h22 == _GEN_4559 ? buffer_1_34 : _GEN_1385; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1387 = 2'h1 == read_ptr[1:0] & 6'h23 == _GEN_4559 ? buffer_1_35 : _GEN_1386; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1388 = 2'h1 == read_ptr[1:0] & 6'h24 == _GEN_4559 ? buffer_1_36 : _GEN_1387; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1389 = 2'h1 == read_ptr[1:0] & 6'h25 == _GEN_4559 ? buffer_1_37 : _GEN_1388; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1390 = 2'h1 == read_ptr[1:0] & 6'h26 == _GEN_4559 ? buffer_1_38 : _GEN_1389; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1391 = 2'h1 == read_ptr[1:0] & 6'h27 == _GEN_4559 ? buffer_1_39 : _GEN_1390; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1392 = 2'h1 == read_ptr[1:0] & 6'h28 == _GEN_4559 ? buffer_1_40 : _GEN_1391; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1393 = 2'h1 == read_ptr[1:0] & 6'h29 == _GEN_4559 ? buffer_1_41 : _GEN_1392; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1394 = 2'h1 == read_ptr[1:0] & 6'h2a == _GEN_4559 ? buffer_1_42 : _GEN_1393; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1395 = 2'h1 == read_ptr[1:0] & 6'h2b == _GEN_4559 ? buffer_1_43 : _GEN_1394; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1396 = 2'h1 == read_ptr[1:0] & 6'h2c == _GEN_4559 ? buffer_1_44 : _GEN_1395; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1397 = 2'h1 == read_ptr[1:0] & 6'h2d == _GEN_4559 ? buffer_1_45 : _GEN_1396; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1398 = 2'h1 == read_ptr[1:0] & 6'h2e == _GEN_4559 ? buffer_1_46 : _GEN_1397; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1399 = 2'h1 == read_ptr[1:0] & 6'h2f == _GEN_4559 ? buffer_1_47 : _GEN_1398; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1400 = 2'h1 == read_ptr[1:0] & 6'h30 == _GEN_4559 ? buffer_1_48 : _GEN_1399; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1401 = 2'h1 == read_ptr[1:0] & 6'h31 == _GEN_4559 ? buffer_1_49 : _GEN_1400; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1402 = 2'h1 == read_ptr[1:0] & 6'h32 == _GEN_4559 ? buffer_1_50 : _GEN_1401; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1403 = 2'h1 == read_ptr[1:0] & 6'h33 == _GEN_4559 ? buffer_1_51 : _GEN_1402; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1404 = 2'h1 == read_ptr[1:0] & 6'h34 == _GEN_4559 ? buffer_1_52 : _GEN_1403; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1405 = 2'h1 == read_ptr[1:0] & 6'h35 == _GEN_4559 ? buffer_1_53 : _GEN_1404; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1406 = 2'h1 == read_ptr[1:0] & 6'h36 == _GEN_4559 ? buffer_1_54 : _GEN_1405; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1407 = 2'h1 == read_ptr[1:0] & 6'h37 == _GEN_4559 ? buffer_1_55 : _GEN_1406; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1408 = 2'h1 == read_ptr[1:0] & 6'h38 == _GEN_4559 ? buffer_1_56 : _GEN_1407; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1409 = 2'h1 == read_ptr[1:0] & 6'h39 == _GEN_4559 ? buffer_1_57 : _GEN_1408; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1410 = 2'h1 == read_ptr[1:0] & 6'h3a == _GEN_4559 ? buffer_1_58 : _GEN_1409; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1411 = 2'h1 == read_ptr[1:0] & 6'h3b == _GEN_4559 ? buffer_1_59 : _GEN_1410; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1412 = 2'h1 == read_ptr[1:0] & 6'h3c == _GEN_4559 ? buffer_1_60 : _GEN_1411; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1413 = 2'h1 == read_ptr[1:0] & 6'h3d == _GEN_4559 ? buffer_1_61 : _GEN_1412; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1414 = 2'h1 == read_ptr[1:0] & 6'h3e == _GEN_4559 ? buffer_1_62 : _GEN_1413; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1415 = 2'h1 == read_ptr[1:0] & 6'h3f == _GEN_4559 ? buffer_1_63 : _GEN_1414; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1416 = 2'h2 == read_ptr[1:0] & 5'h0 == _io_out_activate_3_T_4 ? buffer_2_0 : _GEN_1415; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1417 = 2'h2 == read_ptr[1:0] & 5'h1 == _io_out_activate_3_T_4 ? buffer_2_1 : _GEN_1416; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1418 = 2'h2 == read_ptr[1:0] & 5'h2 == _io_out_activate_3_T_4 ? buffer_2_2 : _GEN_1417; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1419 = 2'h2 == read_ptr[1:0] & 5'h3 == _io_out_activate_3_T_4 ? buffer_2_3 : _GEN_1418; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1420 = 2'h2 == read_ptr[1:0] & 5'h4 == _io_out_activate_3_T_4 ? buffer_2_4 : _GEN_1419; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1421 = 2'h2 == read_ptr[1:0] & 5'h5 == _io_out_activate_3_T_4 ? buffer_2_5 : _GEN_1420; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1422 = 2'h2 == read_ptr[1:0] & 5'h6 == _io_out_activate_3_T_4 ? buffer_2_6 : _GEN_1421; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1423 = 2'h2 == read_ptr[1:0] & 5'h7 == _io_out_activate_3_T_4 ? buffer_2_7 : _GEN_1422; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1424 = 2'h2 == read_ptr[1:0] & 5'h8 == _io_out_activate_3_T_4 ? buffer_2_8 : _GEN_1423; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1425 = 2'h2 == read_ptr[1:0] & 5'h9 == _io_out_activate_3_T_4 ? buffer_2_9 : _GEN_1424; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1426 = 2'h2 == read_ptr[1:0] & 5'ha == _io_out_activate_3_T_4 ? buffer_2_10 : _GEN_1425; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1427 = 2'h2 == read_ptr[1:0] & 5'hb == _io_out_activate_3_T_4 ? buffer_2_11 : _GEN_1426; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1428 = 2'h2 == read_ptr[1:0] & 5'hc == _io_out_activate_3_T_4 ? buffer_2_12 : _GEN_1427; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1429 = 2'h2 == read_ptr[1:0] & 5'hd == _io_out_activate_3_T_4 ? buffer_2_13 : _GEN_1428; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1430 = 2'h2 == read_ptr[1:0] & 5'he == _io_out_activate_3_T_4 ? buffer_2_14 : _GEN_1429; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1431 = 2'h2 == read_ptr[1:0] & 5'hf == _io_out_activate_3_T_4 ? buffer_2_15 : _GEN_1430; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1432 = 2'h2 == read_ptr[1:0] & 5'h10 == _io_out_activate_3_T_4 ? buffer_2_16 : _GEN_1431; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1433 = 2'h2 == read_ptr[1:0] & 5'h11 == _io_out_activate_3_T_4 ? buffer_2_17 : _GEN_1432; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1434 = 2'h2 == read_ptr[1:0] & 5'h12 == _io_out_activate_3_T_4 ? buffer_2_18 : _GEN_1433; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1435 = 2'h2 == read_ptr[1:0] & 5'h13 == _io_out_activate_3_T_4 ? buffer_2_19 : _GEN_1434; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1436 = 2'h2 == read_ptr[1:0] & 5'h14 == _io_out_activate_3_T_4 ? buffer_2_20 : _GEN_1435; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1437 = 2'h2 == read_ptr[1:0] & 5'h15 == _io_out_activate_3_T_4 ? buffer_2_21 : _GEN_1436; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1438 = 2'h2 == read_ptr[1:0] & 5'h16 == _io_out_activate_3_T_4 ? buffer_2_22 : _GEN_1437; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1439 = 2'h2 == read_ptr[1:0] & 5'h17 == _io_out_activate_3_T_4 ? buffer_2_23 : _GEN_1438; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1440 = 2'h2 == read_ptr[1:0] & 5'h18 == _io_out_activate_3_T_4 ? buffer_2_24 : _GEN_1439; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1441 = 2'h2 == read_ptr[1:0] & 5'h19 == _io_out_activate_3_T_4 ? buffer_2_25 : _GEN_1440; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1442 = 2'h2 == read_ptr[1:0] & 5'h1a == _io_out_activate_3_T_4 ? buffer_2_26 : _GEN_1441; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1443 = 2'h2 == read_ptr[1:0] & 5'h1b == _io_out_activate_3_T_4 ? buffer_2_27 : _GEN_1442; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1444 = 2'h2 == read_ptr[1:0] & 5'h1c == _io_out_activate_3_T_4 ? buffer_2_28 : _GEN_1443; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1445 = 2'h2 == read_ptr[1:0] & 5'h1d == _io_out_activate_3_T_4 ? buffer_2_29 : _GEN_1444; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1446 = 2'h2 == read_ptr[1:0] & 5'h1e == _io_out_activate_3_T_4 ? buffer_2_30 : _GEN_1445; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1447 = 2'h2 == read_ptr[1:0] & 5'h1f == _io_out_activate_3_T_4 ? buffer_2_31 : _GEN_1446; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1448 = 2'h2 == read_ptr[1:0] & 6'h20 == _GEN_4559 ? buffer_2_32 : _GEN_1447; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1449 = 2'h2 == read_ptr[1:0] & 6'h21 == _GEN_4559 ? buffer_2_33 : _GEN_1448; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1450 = 2'h2 == read_ptr[1:0] & 6'h22 == _GEN_4559 ? buffer_2_34 : _GEN_1449; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1451 = 2'h2 == read_ptr[1:0] & 6'h23 == _GEN_4559 ? buffer_2_35 : _GEN_1450; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1452 = 2'h2 == read_ptr[1:0] & 6'h24 == _GEN_4559 ? buffer_2_36 : _GEN_1451; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1453 = 2'h2 == read_ptr[1:0] & 6'h25 == _GEN_4559 ? buffer_2_37 : _GEN_1452; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1454 = 2'h2 == read_ptr[1:0] & 6'h26 == _GEN_4559 ? buffer_2_38 : _GEN_1453; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1455 = 2'h2 == read_ptr[1:0] & 6'h27 == _GEN_4559 ? buffer_2_39 : _GEN_1454; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1456 = 2'h2 == read_ptr[1:0] & 6'h28 == _GEN_4559 ? buffer_2_40 : _GEN_1455; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1457 = 2'h2 == read_ptr[1:0] & 6'h29 == _GEN_4559 ? buffer_2_41 : _GEN_1456; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1458 = 2'h2 == read_ptr[1:0] & 6'h2a == _GEN_4559 ? buffer_2_42 : _GEN_1457; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1459 = 2'h2 == read_ptr[1:0] & 6'h2b == _GEN_4559 ? buffer_2_43 : _GEN_1458; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1460 = 2'h2 == read_ptr[1:0] & 6'h2c == _GEN_4559 ? buffer_2_44 : _GEN_1459; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1461 = 2'h2 == read_ptr[1:0] & 6'h2d == _GEN_4559 ? buffer_2_45 : _GEN_1460; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1462 = 2'h2 == read_ptr[1:0] & 6'h2e == _GEN_4559 ? buffer_2_46 : _GEN_1461; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1463 = 2'h2 == read_ptr[1:0] & 6'h2f == _GEN_4559 ? buffer_2_47 : _GEN_1462; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1464 = 2'h2 == read_ptr[1:0] & 6'h30 == _GEN_4559 ? buffer_2_48 : _GEN_1463; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1465 = 2'h2 == read_ptr[1:0] & 6'h31 == _GEN_4559 ? buffer_2_49 : _GEN_1464; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1466 = 2'h2 == read_ptr[1:0] & 6'h32 == _GEN_4559 ? buffer_2_50 : _GEN_1465; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1467 = 2'h2 == read_ptr[1:0] & 6'h33 == _GEN_4559 ? buffer_2_51 : _GEN_1466; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1468 = 2'h2 == read_ptr[1:0] & 6'h34 == _GEN_4559 ? buffer_2_52 : _GEN_1467; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1469 = 2'h2 == read_ptr[1:0] & 6'h35 == _GEN_4559 ? buffer_2_53 : _GEN_1468; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1470 = 2'h2 == read_ptr[1:0] & 6'h36 == _GEN_4559 ? buffer_2_54 : _GEN_1469; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1471 = 2'h2 == read_ptr[1:0] & 6'h37 == _GEN_4559 ? buffer_2_55 : _GEN_1470; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1472 = 2'h2 == read_ptr[1:0] & 6'h38 == _GEN_4559 ? buffer_2_56 : _GEN_1471; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1473 = 2'h2 == read_ptr[1:0] & 6'h39 == _GEN_4559 ? buffer_2_57 : _GEN_1472; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1474 = 2'h2 == read_ptr[1:0] & 6'h3a == _GEN_4559 ? buffer_2_58 : _GEN_1473; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1475 = 2'h2 == read_ptr[1:0] & 6'h3b == _GEN_4559 ? buffer_2_59 : _GEN_1474; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1476 = 2'h2 == read_ptr[1:0] & 6'h3c == _GEN_4559 ? buffer_2_60 : _GEN_1475; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1477 = 2'h2 == read_ptr[1:0] & 6'h3d == _GEN_4559 ? buffer_2_61 : _GEN_1476; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1478 = 2'h2 == read_ptr[1:0] & 6'h3e == _GEN_4559 ? buffer_2_62 : _GEN_1477; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1479 = 2'h2 == read_ptr[1:0] & 6'h3f == _GEN_4559 ? buffer_2_63 : _GEN_1478; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1480 = 2'h3 == read_ptr[1:0] & 5'h0 == _io_out_activate_3_T_4 ? buffer_3_0 : _GEN_1479; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1481 = 2'h3 == read_ptr[1:0] & 5'h1 == _io_out_activate_3_T_4 ? buffer_3_1 : _GEN_1480; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1482 = 2'h3 == read_ptr[1:0] & 5'h2 == _io_out_activate_3_T_4 ? buffer_3_2 : _GEN_1481; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1483 = 2'h3 == read_ptr[1:0] & 5'h3 == _io_out_activate_3_T_4 ? buffer_3_3 : _GEN_1482; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1484 = 2'h3 == read_ptr[1:0] & 5'h4 == _io_out_activate_3_T_4 ? buffer_3_4 : _GEN_1483; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1485 = 2'h3 == read_ptr[1:0] & 5'h5 == _io_out_activate_3_T_4 ? buffer_3_5 : _GEN_1484; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1486 = 2'h3 == read_ptr[1:0] & 5'h6 == _io_out_activate_3_T_4 ? buffer_3_6 : _GEN_1485; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1487 = 2'h3 == read_ptr[1:0] & 5'h7 == _io_out_activate_3_T_4 ? buffer_3_7 : _GEN_1486; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1488 = 2'h3 == read_ptr[1:0] & 5'h8 == _io_out_activate_3_T_4 ? buffer_3_8 : _GEN_1487; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1489 = 2'h3 == read_ptr[1:0] & 5'h9 == _io_out_activate_3_T_4 ? buffer_3_9 : _GEN_1488; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1490 = 2'h3 == read_ptr[1:0] & 5'ha == _io_out_activate_3_T_4 ? buffer_3_10 : _GEN_1489; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1491 = 2'h3 == read_ptr[1:0] & 5'hb == _io_out_activate_3_T_4 ? buffer_3_11 : _GEN_1490; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1492 = 2'h3 == read_ptr[1:0] & 5'hc == _io_out_activate_3_T_4 ? buffer_3_12 : _GEN_1491; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1493 = 2'h3 == read_ptr[1:0] & 5'hd == _io_out_activate_3_T_4 ? buffer_3_13 : _GEN_1492; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1494 = 2'h3 == read_ptr[1:0] & 5'he == _io_out_activate_3_T_4 ? buffer_3_14 : _GEN_1493; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1495 = 2'h3 == read_ptr[1:0] & 5'hf == _io_out_activate_3_T_4 ? buffer_3_15 : _GEN_1494; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1496 = 2'h3 == read_ptr[1:0] & 5'h10 == _io_out_activate_3_T_4 ? buffer_3_16 : _GEN_1495; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1497 = 2'h3 == read_ptr[1:0] & 5'h11 == _io_out_activate_3_T_4 ? buffer_3_17 : _GEN_1496; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1498 = 2'h3 == read_ptr[1:0] & 5'h12 == _io_out_activate_3_T_4 ? buffer_3_18 : _GEN_1497; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1499 = 2'h3 == read_ptr[1:0] & 5'h13 == _io_out_activate_3_T_4 ? buffer_3_19 : _GEN_1498; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1500 = 2'h3 == read_ptr[1:0] & 5'h14 == _io_out_activate_3_T_4 ? buffer_3_20 : _GEN_1499; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1501 = 2'h3 == read_ptr[1:0] & 5'h15 == _io_out_activate_3_T_4 ? buffer_3_21 : _GEN_1500; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1502 = 2'h3 == read_ptr[1:0] & 5'h16 == _io_out_activate_3_T_4 ? buffer_3_22 : _GEN_1501; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1503 = 2'h3 == read_ptr[1:0] & 5'h17 == _io_out_activate_3_T_4 ? buffer_3_23 : _GEN_1502; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1504 = 2'h3 == read_ptr[1:0] & 5'h18 == _io_out_activate_3_T_4 ? buffer_3_24 : _GEN_1503; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1505 = 2'h3 == read_ptr[1:0] & 5'h19 == _io_out_activate_3_T_4 ? buffer_3_25 : _GEN_1504; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1506 = 2'h3 == read_ptr[1:0] & 5'h1a == _io_out_activate_3_T_4 ? buffer_3_26 : _GEN_1505; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1507 = 2'h3 == read_ptr[1:0] & 5'h1b == _io_out_activate_3_T_4 ? buffer_3_27 : _GEN_1506; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1508 = 2'h3 == read_ptr[1:0] & 5'h1c == _io_out_activate_3_T_4 ? buffer_3_28 : _GEN_1507; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1509 = 2'h3 == read_ptr[1:0] & 5'h1d == _io_out_activate_3_T_4 ? buffer_3_29 : _GEN_1508; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1510 = 2'h3 == read_ptr[1:0] & 5'h1e == _io_out_activate_3_T_4 ? buffer_3_30 : _GEN_1509; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1511 = 2'h3 == read_ptr[1:0] & 5'h1f == _io_out_activate_3_T_4 ? buffer_3_31 : _GEN_1510; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1512 = 2'h3 == read_ptr[1:0] & 6'h20 == _GEN_4559 ? buffer_3_32 : _GEN_1511; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1513 = 2'h3 == read_ptr[1:0] & 6'h21 == _GEN_4559 ? buffer_3_33 : _GEN_1512; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1514 = 2'h3 == read_ptr[1:0] & 6'h22 == _GEN_4559 ? buffer_3_34 : _GEN_1513; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1515 = 2'h3 == read_ptr[1:0] & 6'h23 == _GEN_4559 ? buffer_3_35 : _GEN_1514; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1516 = 2'h3 == read_ptr[1:0] & 6'h24 == _GEN_4559 ? buffer_3_36 : _GEN_1515; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1517 = 2'h3 == read_ptr[1:0] & 6'h25 == _GEN_4559 ? buffer_3_37 : _GEN_1516; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1518 = 2'h3 == read_ptr[1:0] & 6'h26 == _GEN_4559 ? buffer_3_38 : _GEN_1517; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1519 = 2'h3 == read_ptr[1:0] & 6'h27 == _GEN_4559 ? buffer_3_39 : _GEN_1518; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1520 = 2'h3 == read_ptr[1:0] & 6'h28 == _GEN_4559 ? buffer_3_40 : _GEN_1519; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1521 = 2'h3 == read_ptr[1:0] & 6'h29 == _GEN_4559 ? buffer_3_41 : _GEN_1520; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1522 = 2'h3 == read_ptr[1:0] & 6'h2a == _GEN_4559 ? buffer_3_42 : _GEN_1521; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1523 = 2'h3 == read_ptr[1:0] & 6'h2b == _GEN_4559 ? buffer_3_43 : _GEN_1522; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1524 = 2'h3 == read_ptr[1:0] & 6'h2c == _GEN_4559 ? buffer_3_44 : _GEN_1523; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1525 = 2'h3 == read_ptr[1:0] & 6'h2d == _GEN_4559 ? buffer_3_45 : _GEN_1524; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1526 = 2'h3 == read_ptr[1:0] & 6'h2e == _GEN_4559 ? buffer_3_46 : _GEN_1525; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1527 = 2'h3 == read_ptr[1:0] & 6'h2f == _GEN_4559 ? buffer_3_47 : _GEN_1526; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1528 = 2'h3 == read_ptr[1:0] & 6'h30 == _GEN_4559 ? buffer_3_48 : _GEN_1527; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1529 = 2'h3 == read_ptr[1:0] & 6'h31 == _GEN_4559 ? buffer_3_49 : _GEN_1528; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1530 = 2'h3 == read_ptr[1:0] & 6'h32 == _GEN_4559 ? buffer_3_50 : _GEN_1529; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1531 = 2'h3 == read_ptr[1:0] & 6'h33 == _GEN_4559 ? buffer_3_51 : _GEN_1530; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1532 = 2'h3 == read_ptr[1:0] & 6'h34 == _GEN_4559 ? buffer_3_52 : _GEN_1531; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1533 = 2'h3 == read_ptr[1:0] & 6'h35 == _GEN_4559 ? buffer_3_53 : _GEN_1532; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1534 = 2'h3 == read_ptr[1:0] & 6'h36 == _GEN_4559 ? buffer_3_54 : _GEN_1533; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1535 = 2'h3 == read_ptr[1:0] & 6'h37 == _GEN_4559 ? buffer_3_55 : _GEN_1534; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1536 = 2'h3 == read_ptr[1:0] & 6'h38 == _GEN_4559 ? buffer_3_56 : _GEN_1535; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1537 = 2'h3 == read_ptr[1:0] & 6'h39 == _GEN_4559 ? buffer_3_57 : _GEN_1536; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1538 = 2'h3 == read_ptr[1:0] & 6'h3a == _GEN_4559 ? buffer_3_58 : _GEN_1537; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1539 = 2'h3 == read_ptr[1:0] & 6'h3b == _GEN_4559 ? buffer_3_59 : _GEN_1538; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1540 = 2'h3 == read_ptr[1:0] & 6'h3c == _GEN_4559 ? buffer_3_60 : _GEN_1539; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1541 = 2'h3 == read_ptr[1:0] & 6'h3d == _GEN_4559 ? buffer_3_61 : _GEN_1540; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1542 = 2'h3 == read_ptr[1:0] & 6'h3e == _GEN_4559 ? buffer_3_62 : _GEN_1541; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1543 = 2'h3 == read_ptr[1:0] & 6'h3f == _GEN_4559 ? buffer_3_63 : _GEN_1542; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1544 = 5'h3 < flow_ptr & flow_ptr <= 5'hb ? _GEN_1543 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [5:0] _io_out_activate_4_T_2 = 6'h20 + _io_out_activate_0_T_1; // @[Activation_Buffer.scala 76:88]
  wire [5:0] _io_out_activate_4_T_4 = _io_out_activate_4_T_2 - 6'h5; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_1546 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_activate_4_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1547 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_activate_4_T_4 ? buffer_0_2 : _GEN_1546; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1548 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_activate_4_T_4 ? buffer_0_3 : _GEN_1547; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1549 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_activate_4_T_4 ? buffer_0_4 : _GEN_1548; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1550 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_activate_4_T_4 ? buffer_0_5 : _GEN_1549; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1551 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_activate_4_T_4 ? buffer_0_6 : _GEN_1550; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1552 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_activate_4_T_4 ? buffer_0_7 : _GEN_1551; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1553 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_activate_4_T_4 ? buffer_0_8 : _GEN_1552; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1554 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_activate_4_T_4 ? buffer_0_9 : _GEN_1553; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1555 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_activate_4_T_4 ? buffer_0_10 : _GEN_1554; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1556 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_activate_4_T_4 ? buffer_0_11 : _GEN_1555; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1557 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_activate_4_T_4 ? buffer_0_12 : _GEN_1556; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1558 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_activate_4_T_4 ? buffer_0_13 : _GEN_1557; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1559 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_activate_4_T_4 ? buffer_0_14 : _GEN_1558; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1560 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_activate_4_T_4 ? buffer_0_15 : _GEN_1559; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1561 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_activate_4_T_4 ? buffer_0_16 : _GEN_1560; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1562 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_activate_4_T_4 ? buffer_0_17 : _GEN_1561; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1563 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_activate_4_T_4 ? buffer_0_18 : _GEN_1562; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1564 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_activate_4_T_4 ? buffer_0_19 : _GEN_1563; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1565 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_activate_4_T_4 ? buffer_0_20 : _GEN_1564; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1566 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_activate_4_T_4 ? buffer_0_21 : _GEN_1565; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1567 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_activate_4_T_4 ? buffer_0_22 : _GEN_1566; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1568 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_activate_4_T_4 ? buffer_0_23 : _GEN_1567; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1569 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_activate_4_T_4 ? buffer_0_24 : _GEN_1568; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1570 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_activate_4_T_4 ? buffer_0_25 : _GEN_1569; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1571 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_activate_4_T_4 ? buffer_0_26 : _GEN_1570; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1572 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_activate_4_T_4 ? buffer_0_27 : _GEN_1571; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1573 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_activate_4_T_4 ? buffer_0_28 : _GEN_1572; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1574 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_activate_4_T_4 ? buffer_0_29 : _GEN_1573; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1575 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_activate_4_T_4 ? buffer_0_30 : _GEN_1574; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1576 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_activate_4_T_4 ? buffer_0_31 : _GEN_1575; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1577 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_activate_4_T_4 ? buffer_0_32 : _GEN_1576; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1578 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_activate_4_T_4 ? buffer_0_33 : _GEN_1577; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1579 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_activate_4_T_4 ? buffer_0_34 : _GEN_1578; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1580 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_activate_4_T_4 ? buffer_0_35 : _GEN_1579; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1581 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_activate_4_T_4 ? buffer_0_36 : _GEN_1580; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1582 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_activate_4_T_4 ? buffer_0_37 : _GEN_1581; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1583 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_activate_4_T_4 ? buffer_0_38 : _GEN_1582; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1584 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_activate_4_T_4 ? buffer_0_39 : _GEN_1583; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1585 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_activate_4_T_4 ? buffer_0_40 : _GEN_1584; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1586 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_activate_4_T_4 ? buffer_0_41 : _GEN_1585; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1587 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_activate_4_T_4 ? buffer_0_42 : _GEN_1586; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1588 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_activate_4_T_4 ? buffer_0_43 : _GEN_1587; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1589 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_activate_4_T_4 ? buffer_0_44 : _GEN_1588; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1590 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_activate_4_T_4 ? buffer_0_45 : _GEN_1589; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1591 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_activate_4_T_4 ? buffer_0_46 : _GEN_1590; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1592 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_activate_4_T_4 ? buffer_0_47 : _GEN_1591; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1593 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_activate_4_T_4 ? buffer_0_48 : _GEN_1592; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1594 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_activate_4_T_4 ? buffer_0_49 : _GEN_1593; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1595 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_activate_4_T_4 ? buffer_0_50 : _GEN_1594; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1596 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_activate_4_T_4 ? buffer_0_51 : _GEN_1595; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1597 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_activate_4_T_4 ? buffer_0_52 : _GEN_1596; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1598 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_activate_4_T_4 ? buffer_0_53 : _GEN_1597; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1599 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_activate_4_T_4 ? buffer_0_54 : _GEN_1598; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1600 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_activate_4_T_4 ? buffer_0_55 : _GEN_1599; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1601 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_activate_4_T_4 ? buffer_0_56 : _GEN_1600; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1602 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_activate_4_T_4 ? buffer_0_57 : _GEN_1601; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1603 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_activate_4_T_4 ? buffer_0_58 : _GEN_1602; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1604 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_activate_4_T_4 ? buffer_0_59 : _GEN_1603; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1605 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_activate_4_T_4 ? buffer_0_60 : _GEN_1604; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1606 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_activate_4_T_4 ? buffer_0_61 : _GEN_1605; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1607 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_activate_4_T_4 ? buffer_0_62 : _GEN_1606; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1608 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_activate_4_T_4 ? buffer_0_63 : _GEN_1607; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1609 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_activate_4_T_4 ? buffer_1_0 : _GEN_1608; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1610 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_activate_4_T_4 ? buffer_1_1 : _GEN_1609; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1611 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_activate_4_T_4 ? buffer_1_2 : _GEN_1610; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1612 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_activate_4_T_4 ? buffer_1_3 : _GEN_1611; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1613 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_activate_4_T_4 ? buffer_1_4 : _GEN_1612; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1614 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_activate_4_T_4 ? buffer_1_5 : _GEN_1613; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1615 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_activate_4_T_4 ? buffer_1_6 : _GEN_1614; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1616 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_activate_4_T_4 ? buffer_1_7 : _GEN_1615; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1617 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_activate_4_T_4 ? buffer_1_8 : _GEN_1616; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1618 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_activate_4_T_4 ? buffer_1_9 : _GEN_1617; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1619 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_activate_4_T_4 ? buffer_1_10 : _GEN_1618; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1620 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_activate_4_T_4 ? buffer_1_11 : _GEN_1619; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1621 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_activate_4_T_4 ? buffer_1_12 : _GEN_1620; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1622 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_activate_4_T_4 ? buffer_1_13 : _GEN_1621; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1623 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_activate_4_T_4 ? buffer_1_14 : _GEN_1622; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1624 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_activate_4_T_4 ? buffer_1_15 : _GEN_1623; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1625 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_activate_4_T_4 ? buffer_1_16 : _GEN_1624; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1626 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_activate_4_T_4 ? buffer_1_17 : _GEN_1625; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1627 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_activate_4_T_4 ? buffer_1_18 : _GEN_1626; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1628 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_activate_4_T_4 ? buffer_1_19 : _GEN_1627; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1629 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_activate_4_T_4 ? buffer_1_20 : _GEN_1628; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1630 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_activate_4_T_4 ? buffer_1_21 : _GEN_1629; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1631 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_activate_4_T_4 ? buffer_1_22 : _GEN_1630; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1632 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_activate_4_T_4 ? buffer_1_23 : _GEN_1631; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1633 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_activate_4_T_4 ? buffer_1_24 : _GEN_1632; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1634 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_activate_4_T_4 ? buffer_1_25 : _GEN_1633; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1635 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_activate_4_T_4 ? buffer_1_26 : _GEN_1634; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1636 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_activate_4_T_4 ? buffer_1_27 : _GEN_1635; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1637 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_activate_4_T_4 ? buffer_1_28 : _GEN_1636; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1638 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_activate_4_T_4 ? buffer_1_29 : _GEN_1637; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1639 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_activate_4_T_4 ? buffer_1_30 : _GEN_1638; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1640 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_activate_4_T_4 ? buffer_1_31 : _GEN_1639; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1641 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_activate_4_T_4 ? buffer_1_32 : _GEN_1640; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1642 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_activate_4_T_4 ? buffer_1_33 : _GEN_1641; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1643 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_activate_4_T_4 ? buffer_1_34 : _GEN_1642; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1644 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_activate_4_T_4 ? buffer_1_35 : _GEN_1643; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1645 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_activate_4_T_4 ? buffer_1_36 : _GEN_1644; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1646 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_activate_4_T_4 ? buffer_1_37 : _GEN_1645; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1647 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_activate_4_T_4 ? buffer_1_38 : _GEN_1646; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1648 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_activate_4_T_4 ? buffer_1_39 : _GEN_1647; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1649 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_activate_4_T_4 ? buffer_1_40 : _GEN_1648; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1650 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_activate_4_T_4 ? buffer_1_41 : _GEN_1649; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1651 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_activate_4_T_4 ? buffer_1_42 : _GEN_1650; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1652 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_activate_4_T_4 ? buffer_1_43 : _GEN_1651; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1653 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_activate_4_T_4 ? buffer_1_44 : _GEN_1652; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1654 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_activate_4_T_4 ? buffer_1_45 : _GEN_1653; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1655 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_activate_4_T_4 ? buffer_1_46 : _GEN_1654; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1656 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_activate_4_T_4 ? buffer_1_47 : _GEN_1655; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1657 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_activate_4_T_4 ? buffer_1_48 : _GEN_1656; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1658 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_activate_4_T_4 ? buffer_1_49 : _GEN_1657; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1659 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_activate_4_T_4 ? buffer_1_50 : _GEN_1658; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1660 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_activate_4_T_4 ? buffer_1_51 : _GEN_1659; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1661 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_activate_4_T_4 ? buffer_1_52 : _GEN_1660; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1662 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_activate_4_T_4 ? buffer_1_53 : _GEN_1661; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1663 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_activate_4_T_4 ? buffer_1_54 : _GEN_1662; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1664 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_activate_4_T_4 ? buffer_1_55 : _GEN_1663; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1665 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_activate_4_T_4 ? buffer_1_56 : _GEN_1664; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1666 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_activate_4_T_4 ? buffer_1_57 : _GEN_1665; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1667 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_activate_4_T_4 ? buffer_1_58 : _GEN_1666; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1668 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_activate_4_T_4 ? buffer_1_59 : _GEN_1667; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1669 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_activate_4_T_4 ? buffer_1_60 : _GEN_1668; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1670 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_activate_4_T_4 ? buffer_1_61 : _GEN_1669; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1671 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_activate_4_T_4 ? buffer_1_62 : _GEN_1670; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1672 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_activate_4_T_4 ? buffer_1_63 : _GEN_1671; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1673 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_activate_4_T_4 ? buffer_2_0 : _GEN_1672; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1674 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_activate_4_T_4 ? buffer_2_1 : _GEN_1673; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1675 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_activate_4_T_4 ? buffer_2_2 : _GEN_1674; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1676 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_activate_4_T_4 ? buffer_2_3 : _GEN_1675; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1677 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_activate_4_T_4 ? buffer_2_4 : _GEN_1676; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1678 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_activate_4_T_4 ? buffer_2_5 : _GEN_1677; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1679 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_activate_4_T_4 ? buffer_2_6 : _GEN_1678; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1680 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_activate_4_T_4 ? buffer_2_7 : _GEN_1679; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1681 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_activate_4_T_4 ? buffer_2_8 : _GEN_1680; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1682 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_activate_4_T_4 ? buffer_2_9 : _GEN_1681; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1683 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_activate_4_T_4 ? buffer_2_10 : _GEN_1682; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1684 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_activate_4_T_4 ? buffer_2_11 : _GEN_1683; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1685 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_activate_4_T_4 ? buffer_2_12 : _GEN_1684; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1686 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_activate_4_T_4 ? buffer_2_13 : _GEN_1685; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1687 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_activate_4_T_4 ? buffer_2_14 : _GEN_1686; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1688 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_activate_4_T_4 ? buffer_2_15 : _GEN_1687; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1689 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_activate_4_T_4 ? buffer_2_16 : _GEN_1688; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1690 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_activate_4_T_4 ? buffer_2_17 : _GEN_1689; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1691 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_activate_4_T_4 ? buffer_2_18 : _GEN_1690; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1692 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_activate_4_T_4 ? buffer_2_19 : _GEN_1691; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1693 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_activate_4_T_4 ? buffer_2_20 : _GEN_1692; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1694 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_activate_4_T_4 ? buffer_2_21 : _GEN_1693; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1695 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_activate_4_T_4 ? buffer_2_22 : _GEN_1694; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1696 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_activate_4_T_4 ? buffer_2_23 : _GEN_1695; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1697 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_activate_4_T_4 ? buffer_2_24 : _GEN_1696; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1698 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_activate_4_T_4 ? buffer_2_25 : _GEN_1697; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1699 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_activate_4_T_4 ? buffer_2_26 : _GEN_1698; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1700 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_activate_4_T_4 ? buffer_2_27 : _GEN_1699; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1701 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_activate_4_T_4 ? buffer_2_28 : _GEN_1700; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1702 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_activate_4_T_4 ? buffer_2_29 : _GEN_1701; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1703 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_activate_4_T_4 ? buffer_2_30 : _GEN_1702; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1704 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_activate_4_T_4 ? buffer_2_31 : _GEN_1703; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1705 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_activate_4_T_4 ? buffer_2_32 : _GEN_1704; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1706 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_activate_4_T_4 ? buffer_2_33 : _GEN_1705; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1707 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_activate_4_T_4 ? buffer_2_34 : _GEN_1706; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1708 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_activate_4_T_4 ? buffer_2_35 : _GEN_1707; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1709 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_activate_4_T_4 ? buffer_2_36 : _GEN_1708; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1710 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_activate_4_T_4 ? buffer_2_37 : _GEN_1709; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1711 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_activate_4_T_4 ? buffer_2_38 : _GEN_1710; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1712 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_activate_4_T_4 ? buffer_2_39 : _GEN_1711; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1713 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_activate_4_T_4 ? buffer_2_40 : _GEN_1712; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1714 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_activate_4_T_4 ? buffer_2_41 : _GEN_1713; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1715 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_activate_4_T_4 ? buffer_2_42 : _GEN_1714; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1716 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_activate_4_T_4 ? buffer_2_43 : _GEN_1715; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1717 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_activate_4_T_4 ? buffer_2_44 : _GEN_1716; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1718 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_activate_4_T_4 ? buffer_2_45 : _GEN_1717; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1719 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_activate_4_T_4 ? buffer_2_46 : _GEN_1718; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1720 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_activate_4_T_4 ? buffer_2_47 : _GEN_1719; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1721 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_activate_4_T_4 ? buffer_2_48 : _GEN_1720; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1722 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_activate_4_T_4 ? buffer_2_49 : _GEN_1721; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1723 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_activate_4_T_4 ? buffer_2_50 : _GEN_1722; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1724 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_activate_4_T_4 ? buffer_2_51 : _GEN_1723; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1725 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_activate_4_T_4 ? buffer_2_52 : _GEN_1724; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1726 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_activate_4_T_4 ? buffer_2_53 : _GEN_1725; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1727 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_activate_4_T_4 ? buffer_2_54 : _GEN_1726; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1728 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_activate_4_T_4 ? buffer_2_55 : _GEN_1727; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1729 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_activate_4_T_4 ? buffer_2_56 : _GEN_1728; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1730 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_activate_4_T_4 ? buffer_2_57 : _GEN_1729; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1731 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_activate_4_T_4 ? buffer_2_58 : _GEN_1730; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1732 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_activate_4_T_4 ? buffer_2_59 : _GEN_1731; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1733 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_activate_4_T_4 ? buffer_2_60 : _GEN_1732; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1734 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_activate_4_T_4 ? buffer_2_61 : _GEN_1733; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1735 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_activate_4_T_4 ? buffer_2_62 : _GEN_1734; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1736 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_activate_4_T_4 ? buffer_2_63 : _GEN_1735; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1737 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_activate_4_T_4 ? buffer_3_0 : _GEN_1736; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1738 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_activate_4_T_4 ? buffer_3_1 : _GEN_1737; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1739 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_activate_4_T_4 ? buffer_3_2 : _GEN_1738; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1740 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_activate_4_T_4 ? buffer_3_3 : _GEN_1739; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1741 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_activate_4_T_4 ? buffer_3_4 : _GEN_1740; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1742 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_activate_4_T_4 ? buffer_3_5 : _GEN_1741; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1743 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_activate_4_T_4 ? buffer_3_6 : _GEN_1742; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1744 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_activate_4_T_4 ? buffer_3_7 : _GEN_1743; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1745 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_activate_4_T_4 ? buffer_3_8 : _GEN_1744; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1746 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_activate_4_T_4 ? buffer_3_9 : _GEN_1745; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1747 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_activate_4_T_4 ? buffer_3_10 : _GEN_1746; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1748 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_activate_4_T_4 ? buffer_3_11 : _GEN_1747; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1749 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_activate_4_T_4 ? buffer_3_12 : _GEN_1748; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1750 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_activate_4_T_4 ? buffer_3_13 : _GEN_1749; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1751 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_activate_4_T_4 ? buffer_3_14 : _GEN_1750; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1752 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_activate_4_T_4 ? buffer_3_15 : _GEN_1751; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1753 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_activate_4_T_4 ? buffer_3_16 : _GEN_1752; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1754 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_activate_4_T_4 ? buffer_3_17 : _GEN_1753; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1755 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_activate_4_T_4 ? buffer_3_18 : _GEN_1754; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1756 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_activate_4_T_4 ? buffer_3_19 : _GEN_1755; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1757 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_activate_4_T_4 ? buffer_3_20 : _GEN_1756; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1758 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_activate_4_T_4 ? buffer_3_21 : _GEN_1757; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1759 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_activate_4_T_4 ? buffer_3_22 : _GEN_1758; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1760 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_activate_4_T_4 ? buffer_3_23 : _GEN_1759; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1761 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_activate_4_T_4 ? buffer_3_24 : _GEN_1760; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1762 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_activate_4_T_4 ? buffer_3_25 : _GEN_1761; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1763 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_activate_4_T_4 ? buffer_3_26 : _GEN_1762; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1764 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_activate_4_T_4 ? buffer_3_27 : _GEN_1763; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1765 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_activate_4_T_4 ? buffer_3_28 : _GEN_1764; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1766 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_activate_4_T_4 ? buffer_3_29 : _GEN_1765; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1767 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_activate_4_T_4 ? buffer_3_30 : _GEN_1766; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1768 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_activate_4_T_4 ? buffer_3_31 : _GEN_1767; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1769 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_activate_4_T_4 ? buffer_3_32 : _GEN_1768; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1770 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_activate_4_T_4 ? buffer_3_33 : _GEN_1769; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1771 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_activate_4_T_4 ? buffer_3_34 : _GEN_1770; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1772 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_activate_4_T_4 ? buffer_3_35 : _GEN_1771; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1773 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_activate_4_T_4 ? buffer_3_36 : _GEN_1772; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1774 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_activate_4_T_4 ? buffer_3_37 : _GEN_1773; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1775 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_activate_4_T_4 ? buffer_3_38 : _GEN_1774; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1776 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_activate_4_T_4 ? buffer_3_39 : _GEN_1775; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1777 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_activate_4_T_4 ? buffer_3_40 : _GEN_1776; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1778 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_activate_4_T_4 ? buffer_3_41 : _GEN_1777; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1779 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_activate_4_T_4 ? buffer_3_42 : _GEN_1778; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1780 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_activate_4_T_4 ? buffer_3_43 : _GEN_1779; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1781 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_activate_4_T_4 ? buffer_3_44 : _GEN_1780; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1782 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_activate_4_T_4 ? buffer_3_45 : _GEN_1781; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1783 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_activate_4_T_4 ? buffer_3_46 : _GEN_1782; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1784 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_activate_4_T_4 ? buffer_3_47 : _GEN_1783; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1785 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_activate_4_T_4 ? buffer_3_48 : _GEN_1784; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1786 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_activate_4_T_4 ? buffer_3_49 : _GEN_1785; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1787 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_activate_4_T_4 ? buffer_3_50 : _GEN_1786; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1788 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_activate_4_T_4 ? buffer_3_51 : _GEN_1787; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1789 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_activate_4_T_4 ? buffer_3_52 : _GEN_1788; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1790 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_activate_4_T_4 ? buffer_3_53 : _GEN_1789; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1791 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_activate_4_T_4 ? buffer_3_54 : _GEN_1790; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1792 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_activate_4_T_4 ? buffer_3_55 : _GEN_1791; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1793 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_activate_4_T_4 ? buffer_3_56 : _GEN_1792; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1794 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_activate_4_T_4 ? buffer_3_57 : _GEN_1793; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1795 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_activate_4_T_4 ? buffer_3_58 : _GEN_1794; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1796 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_activate_4_T_4 ? buffer_3_59 : _GEN_1795; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1797 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_activate_4_T_4 ? buffer_3_60 : _GEN_1796; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1798 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_activate_4_T_4 ? buffer_3_61 : _GEN_1797; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1799 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_activate_4_T_4 ? buffer_3_62 : _GEN_1798; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1800 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_activate_4_T_4 ? buffer_3_63 : _GEN_1799; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1801 = 5'h4 < flow_ptr & flow_ptr <= 5'hc ? _GEN_1800 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [5:0] _io_out_activate_5_T_2 = 6'h28 + _io_out_activate_0_T_1; // @[Activation_Buffer.scala 76:88]
  wire [5:0] _io_out_activate_5_T_4 = _io_out_activate_5_T_2 - 6'h6; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_1803 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_activate_5_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1804 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_activate_5_T_4 ? buffer_0_2 : _GEN_1803; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1805 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_activate_5_T_4 ? buffer_0_3 : _GEN_1804; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1806 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_activate_5_T_4 ? buffer_0_4 : _GEN_1805; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1807 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_activate_5_T_4 ? buffer_0_5 : _GEN_1806; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1808 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_activate_5_T_4 ? buffer_0_6 : _GEN_1807; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1809 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_activate_5_T_4 ? buffer_0_7 : _GEN_1808; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1810 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_activate_5_T_4 ? buffer_0_8 : _GEN_1809; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1811 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_activate_5_T_4 ? buffer_0_9 : _GEN_1810; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1812 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_activate_5_T_4 ? buffer_0_10 : _GEN_1811; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1813 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_activate_5_T_4 ? buffer_0_11 : _GEN_1812; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1814 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_activate_5_T_4 ? buffer_0_12 : _GEN_1813; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1815 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_activate_5_T_4 ? buffer_0_13 : _GEN_1814; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1816 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_activate_5_T_4 ? buffer_0_14 : _GEN_1815; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1817 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_activate_5_T_4 ? buffer_0_15 : _GEN_1816; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1818 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_activate_5_T_4 ? buffer_0_16 : _GEN_1817; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1819 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_activate_5_T_4 ? buffer_0_17 : _GEN_1818; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1820 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_activate_5_T_4 ? buffer_0_18 : _GEN_1819; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1821 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_activate_5_T_4 ? buffer_0_19 : _GEN_1820; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1822 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_activate_5_T_4 ? buffer_0_20 : _GEN_1821; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1823 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_activate_5_T_4 ? buffer_0_21 : _GEN_1822; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1824 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_activate_5_T_4 ? buffer_0_22 : _GEN_1823; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1825 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_activate_5_T_4 ? buffer_0_23 : _GEN_1824; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1826 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_activate_5_T_4 ? buffer_0_24 : _GEN_1825; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1827 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_activate_5_T_4 ? buffer_0_25 : _GEN_1826; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1828 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_activate_5_T_4 ? buffer_0_26 : _GEN_1827; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1829 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_activate_5_T_4 ? buffer_0_27 : _GEN_1828; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1830 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_activate_5_T_4 ? buffer_0_28 : _GEN_1829; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1831 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_activate_5_T_4 ? buffer_0_29 : _GEN_1830; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1832 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_activate_5_T_4 ? buffer_0_30 : _GEN_1831; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1833 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_activate_5_T_4 ? buffer_0_31 : _GEN_1832; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1834 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_activate_5_T_4 ? buffer_0_32 : _GEN_1833; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1835 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_activate_5_T_4 ? buffer_0_33 : _GEN_1834; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1836 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_activate_5_T_4 ? buffer_0_34 : _GEN_1835; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1837 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_activate_5_T_4 ? buffer_0_35 : _GEN_1836; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1838 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_activate_5_T_4 ? buffer_0_36 : _GEN_1837; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1839 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_activate_5_T_4 ? buffer_0_37 : _GEN_1838; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1840 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_activate_5_T_4 ? buffer_0_38 : _GEN_1839; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1841 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_activate_5_T_4 ? buffer_0_39 : _GEN_1840; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1842 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_activate_5_T_4 ? buffer_0_40 : _GEN_1841; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1843 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_activate_5_T_4 ? buffer_0_41 : _GEN_1842; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1844 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_activate_5_T_4 ? buffer_0_42 : _GEN_1843; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1845 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_activate_5_T_4 ? buffer_0_43 : _GEN_1844; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1846 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_activate_5_T_4 ? buffer_0_44 : _GEN_1845; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1847 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_activate_5_T_4 ? buffer_0_45 : _GEN_1846; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1848 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_activate_5_T_4 ? buffer_0_46 : _GEN_1847; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1849 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_activate_5_T_4 ? buffer_0_47 : _GEN_1848; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1850 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_activate_5_T_4 ? buffer_0_48 : _GEN_1849; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1851 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_activate_5_T_4 ? buffer_0_49 : _GEN_1850; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1852 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_activate_5_T_4 ? buffer_0_50 : _GEN_1851; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1853 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_activate_5_T_4 ? buffer_0_51 : _GEN_1852; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1854 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_activate_5_T_4 ? buffer_0_52 : _GEN_1853; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1855 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_activate_5_T_4 ? buffer_0_53 : _GEN_1854; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1856 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_activate_5_T_4 ? buffer_0_54 : _GEN_1855; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1857 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_activate_5_T_4 ? buffer_0_55 : _GEN_1856; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1858 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_activate_5_T_4 ? buffer_0_56 : _GEN_1857; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1859 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_activate_5_T_4 ? buffer_0_57 : _GEN_1858; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1860 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_activate_5_T_4 ? buffer_0_58 : _GEN_1859; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1861 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_activate_5_T_4 ? buffer_0_59 : _GEN_1860; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1862 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_activate_5_T_4 ? buffer_0_60 : _GEN_1861; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1863 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_activate_5_T_4 ? buffer_0_61 : _GEN_1862; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1864 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_activate_5_T_4 ? buffer_0_62 : _GEN_1863; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1865 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_activate_5_T_4 ? buffer_0_63 : _GEN_1864; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1866 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_activate_5_T_4 ? buffer_1_0 : _GEN_1865; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1867 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_activate_5_T_4 ? buffer_1_1 : _GEN_1866; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1868 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_activate_5_T_4 ? buffer_1_2 : _GEN_1867; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1869 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_activate_5_T_4 ? buffer_1_3 : _GEN_1868; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1870 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_activate_5_T_4 ? buffer_1_4 : _GEN_1869; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1871 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_activate_5_T_4 ? buffer_1_5 : _GEN_1870; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1872 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_activate_5_T_4 ? buffer_1_6 : _GEN_1871; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1873 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_activate_5_T_4 ? buffer_1_7 : _GEN_1872; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1874 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_activate_5_T_4 ? buffer_1_8 : _GEN_1873; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1875 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_activate_5_T_4 ? buffer_1_9 : _GEN_1874; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1876 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_activate_5_T_4 ? buffer_1_10 : _GEN_1875; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1877 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_activate_5_T_4 ? buffer_1_11 : _GEN_1876; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1878 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_activate_5_T_4 ? buffer_1_12 : _GEN_1877; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1879 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_activate_5_T_4 ? buffer_1_13 : _GEN_1878; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1880 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_activate_5_T_4 ? buffer_1_14 : _GEN_1879; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1881 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_activate_5_T_4 ? buffer_1_15 : _GEN_1880; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1882 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_activate_5_T_4 ? buffer_1_16 : _GEN_1881; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1883 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_activate_5_T_4 ? buffer_1_17 : _GEN_1882; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1884 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_activate_5_T_4 ? buffer_1_18 : _GEN_1883; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1885 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_activate_5_T_4 ? buffer_1_19 : _GEN_1884; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1886 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_activate_5_T_4 ? buffer_1_20 : _GEN_1885; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1887 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_activate_5_T_4 ? buffer_1_21 : _GEN_1886; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1888 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_activate_5_T_4 ? buffer_1_22 : _GEN_1887; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1889 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_activate_5_T_4 ? buffer_1_23 : _GEN_1888; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1890 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_activate_5_T_4 ? buffer_1_24 : _GEN_1889; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1891 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_activate_5_T_4 ? buffer_1_25 : _GEN_1890; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1892 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_activate_5_T_4 ? buffer_1_26 : _GEN_1891; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1893 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_activate_5_T_4 ? buffer_1_27 : _GEN_1892; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1894 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_activate_5_T_4 ? buffer_1_28 : _GEN_1893; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1895 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_activate_5_T_4 ? buffer_1_29 : _GEN_1894; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1896 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_activate_5_T_4 ? buffer_1_30 : _GEN_1895; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1897 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_activate_5_T_4 ? buffer_1_31 : _GEN_1896; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1898 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_activate_5_T_4 ? buffer_1_32 : _GEN_1897; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1899 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_activate_5_T_4 ? buffer_1_33 : _GEN_1898; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1900 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_activate_5_T_4 ? buffer_1_34 : _GEN_1899; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1901 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_activate_5_T_4 ? buffer_1_35 : _GEN_1900; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1902 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_activate_5_T_4 ? buffer_1_36 : _GEN_1901; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1903 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_activate_5_T_4 ? buffer_1_37 : _GEN_1902; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1904 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_activate_5_T_4 ? buffer_1_38 : _GEN_1903; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1905 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_activate_5_T_4 ? buffer_1_39 : _GEN_1904; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1906 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_activate_5_T_4 ? buffer_1_40 : _GEN_1905; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1907 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_activate_5_T_4 ? buffer_1_41 : _GEN_1906; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1908 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_activate_5_T_4 ? buffer_1_42 : _GEN_1907; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1909 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_activate_5_T_4 ? buffer_1_43 : _GEN_1908; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1910 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_activate_5_T_4 ? buffer_1_44 : _GEN_1909; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1911 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_activate_5_T_4 ? buffer_1_45 : _GEN_1910; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1912 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_activate_5_T_4 ? buffer_1_46 : _GEN_1911; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1913 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_activate_5_T_4 ? buffer_1_47 : _GEN_1912; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1914 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_activate_5_T_4 ? buffer_1_48 : _GEN_1913; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1915 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_activate_5_T_4 ? buffer_1_49 : _GEN_1914; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1916 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_activate_5_T_4 ? buffer_1_50 : _GEN_1915; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1917 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_activate_5_T_4 ? buffer_1_51 : _GEN_1916; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1918 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_activate_5_T_4 ? buffer_1_52 : _GEN_1917; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1919 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_activate_5_T_4 ? buffer_1_53 : _GEN_1918; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1920 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_activate_5_T_4 ? buffer_1_54 : _GEN_1919; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1921 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_activate_5_T_4 ? buffer_1_55 : _GEN_1920; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1922 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_activate_5_T_4 ? buffer_1_56 : _GEN_1921; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1923 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_activate_5_T_4 ? buffer_1_57 : _GEN_1922; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1924 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_activate_5_T_4 ? buffer_1_58 : _GEN_1923; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1925 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_activate_5_T_4 ? buffer_1_59 : _GEN_1924; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1926 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_activate_5_T_4 ? buffer_1_60 : _GEN_1925; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1927 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_activate_5_T_4 ? buffer_1_61 : _GEN_1926; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1928 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_activate_5_T_4 ? buffer_1_62 : _GEN_1927; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1929 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_activate_5_T_4 ? buffer_1_63 : _GEN_1928; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1930 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_activate_5_T_4 ? buffer_2_0 : _GEN_1929; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1931 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_activate_5_T_4 ? buffer_2_1 : _GEN_1930; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1932 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_activate_5_T_4 ? buffer_2_2 : _GEN_1931; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1933 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_activate_5_T_4 ? buffer_2_3 : _GEN_1932; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1934 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_activate_5_T_4 ? buffer_2_4 : _GEN_1933; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1935 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_activate_5_T_4 ? buffer_2_5 : _GEN_1934; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1936 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_activate_5_T_4 ? buffer_2_6 : _GEN_1935; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1937 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_activate_5_T_4 ? buffer_2_7 : _GEN_1936; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1938 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_activate_5_T_4 ? buffer_2_8 : _GEN_1937; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1939 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_activate_5_T_4 ? buffer_2_9 : _GEN_1938; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1940 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_activate_5_T_4 ? buffer_2_10 : _GEN_1939; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1941 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_activate_5_T_4 ? buffer_2_11 : _GEN_1940; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1942 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_activate_5_T_4 ? buffer_2_12 : _GEN_1941; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1943 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_activate_5_T_4 ? buffer_2_13 : _GEN_1942; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1944 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_activate_5_T_4 ? buffer_2_14 : _GEN_1943; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1945 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_activate_5_T_4 ? buffer_2_15 : _GEN_1944; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1946 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_activate_5_T_4 ? buffer_2_16 : _GEN_1945; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1947 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_activate_5_T_4 ? buffer_2_17 : _GEN_1946; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1948 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_activate_5_T_4 ? buffer_2_18 : _GEN_1947; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1949 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_activate_5_T_4 ? buffer_2_19 : _GEN_1948; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1950 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_activate_5_T_4 ? buffer_2_20 : _GEN_1949; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1951 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_activate_5_T_4 ? buffer_2_21 : _GEN_1950; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1952 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_activate_5_T_4 ? buffer_2_22 : _GEN_1951; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1953 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_activate_5_T_4 ? buffer_2_23 : _GEN_1952; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1954 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_activate_5_T_4 ? buffer_2_24 : _GEN_1953; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1955 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_activate_5_T_4 ? buffer_2_25 : _GEN_1954; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1956 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_activate_5_T_4 ? buffer_2_26 : _GEN_1955; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1957 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_activate_5_T_4 ? buffer_2_27 : _GEN_1956; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1958 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_activate_5_T_4 ? buffer_2_28 : _GEN_1957; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1959 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_activate_5_T_4 ? buffer_2_29 : _GEN_1958; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1960 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_activate_5_T_4 ? buffer_2_30 : _GEN_1959; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1961 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_activate_5_T_4 ? buffer_2_31 : _GEN_1960; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1962 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_activate_5_T_4 ? buffer_2_32 : _GEN_1961; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1963 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_activate_5_T_4 ? buffer_2_33 : _GEN_1962; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1964 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_activate_5_T_4 ? buffer_2_34 : _GEN_1963; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1965 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_activate_5_T_4 ? buffer_2_35 : _GEN_1964; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1966 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_activate_5_T_4 ? buffer_2_36 : _GEN_1965; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1967 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_activate_5_T_4 ? buffer_2_37 : _GEN_1966; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1968 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_activate_5_T_4 ? buffer_2_38 : _GEN_1967; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1969 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_activate_5_T_4 ? buffer_2_39 : _GEN_1968; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1970 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_activate_5_T_4 ? buffer_2_40 : _GEN_1969; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1971 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_activate_5_T_4 ? buffer_2_41 : _GEN_1970; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1972 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_activate_5_T_4 ? buffer_2_42 : _GEN_1971; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1973 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_activate_5_T_4 ? buffer_2_43 : _GEN_1972; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1974 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_activate_5_T_4 ? buffer_2_44 : _GEN_1973; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1975 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_activate_5_T_4 ? buffer_2_45 : _GEN_1974; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1976 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_activate_5_T_4 ? buffer_2_46 : _GEN_1975; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1977 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_activate_5_T_4 ? buffer_2_47 : _GEN_1976; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1978 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_activate_5_T_4 ? buffer_2_48 : _GEN_1977; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1979 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_activate_5_T_4 ? buffer_2_49 : _GEN_1978; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1980 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_activate_5_T_4 ? buffer_2_50 : _GEN_1979; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1981 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_activate_5_T_4 ? buffer_2_51 : _GEN_1980; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1982 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_activate_5_T_4 ? buffer_2_52 : _GEN_1981; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1983 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_activate_5_T_4 ? buffer_2_53 : _GEN_1982; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1984 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_activate_5_T_4 ? buffer_2_54 : _GEN_1983; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1985 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_activate_5_T_4 ? buffer_2_55 : _GEN_1984; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1986 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_activate_5_T_4 ? buffer_2_56 : _GEN_1985; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1987 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_activate_5_T_4 ? buffer_2_57 : _GEN_1986; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1988 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_activate_5_T_4 ? buffer_2_58 : _GEN_1987; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1989 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_activate_5_T_4 ? buffer_2_59 : _GEN_1988; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1990 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_activate_5_T_4 ? buffer_2_60 : _GEN_1989; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1991 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_activate_5_T_4 ? buffer_2_61 : _GEN_1990; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1992 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_activate_5_T_4 ? buffer_2_62 : _GEN_1991; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1993 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_activate_5_T_4 ? buffer_2_63 : _GEN_1992; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1994 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_activate_5_T_4 ? buffer_3_0 : _GEN_1993; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1995 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_activate_5_T_4 ? buffer_3_1 : _GEN_1994; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1996 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_activate_5_T_4 ? buffer_3_2 : _GEN_1995; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1997 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_activate_5_T_4 ? buffer_3_3 : _GEN_1996; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1998 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_activate_5_T_4 ? buffer_3_4 : _GEN_1997; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_1999 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_activate_5_T_4 ? buffer_3_5 : _GEN_1998; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2000 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_activate_5_T_4 ? buffer_3_6 : _GEN_1999; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2001 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_activate_5_T_4 ? buffer_3_7 : _GEN_2000; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2002 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_activate_5_T_4 ? buffer_3_8 : _GEN_2001; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2003 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_activate_5_T_4 ? buffer_3_9 : _GEN_2002; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2004 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_activate_5_T_4 ? buffer_3_10 : _GEN_2003; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2005 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_activate_5_T_4 ? buffer_3_11 : _GEN_2004; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2006 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_activate_5_T_4 ? buffer_3_12 : _GEN_2005; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2007 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_activate_5_T_4 ? buffer_3_13 : _GEN_2006; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2008 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_activate_5_T_4 ? buffer_3_14 : _GEN_2007; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2009 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_activate_5_T_4 ? buffer_3_15 : _GEN_2008; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2010 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_activate_5_T_4 ? buffer_3_16 : _GEN_2009; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2011 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_activate_5_T_4 ? buffer_3_17 : _GEN_2010; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2012 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_activate_5_T_4 ? buffer_3_18 : _GEN_2011; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2013 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_activate_5_T_4 ? buffer_3_19 : _GEN_2012; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2014 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_activate_5_T_4 ? buffer_3_20 : _GEN_2013; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2015 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_activate_5_T_4 ? buffer_3_21 : _GEN_2014; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2016 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_activate_5_T_4 ? buffer_3_22 : _GEN_2015; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2017 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_activate_5_T_4 ? buffer_3_23 : _GEN_2016; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2018 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_activate_5_T_4 ? buffer_3_24 : _GEN_2017; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2019 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_activate_5_T_4 ? buffer_3_25 : _GEN_2018; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2020 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_activate_5_T_4 ? buffer_3_26 : _GEN_2019; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2021 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_activate_5_T_4 ? buffer_3_27 : _GEN_2020; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2022 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_activate_5_T_4 ? buffer_3_28 : _GEN_2021; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2023 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_activate_5_T_4 ? buffer_3_29 : _GEN_2022; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2024 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_activate_5_T_4 ? buffer_3_30 : _GEN_2023; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2025 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_activate_5_T_4 ? buffer_3_31 : _GEN_2024; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2026 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_activate_5_T_4 ? buffer_3_32 : _GEN_2025; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2027 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_activate_5_T_4 ? buffer_3_33 : _GEN_2026; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2028 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_activate_5_T_4 ? buffer_3_34 : _GEN_2027; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2029 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_activate_5_T_4 ? buffer_3_35 : _GEN_2028; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2030 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_activate_5_T_4 ? buffer_3_36 : _GEN_2029; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2031 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_activate_5_T_4 ? buffer_3_37 : _GEN_2030; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2032 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_activate_5_T_4 ? buffer_3_38 : _GEN_2031; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2033 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_activate_5_T_4 ? buffer_3_39 : _GEN_2032; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2034 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_activate_5_T_4 ? buffer_3_40 : _GEN_2033; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2035 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_activate_5_T_4 ? buffer_3_41 : _GEN_2034; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2036 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_activate_5_T_4 ? buffer_3_42 : _GEN_2035; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2037 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_activate_5_T_4 ? buffer_3_43 : _GEN_2036; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2038 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_activate_5_T_4 ? buffer_3_44 : _GEN_2037; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2039 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_activate_5_T_4 ? buffer_3_45 : _GEN_2038; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2040 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_activate_5_T_4 ? buffer_3_46 : _GEN_2039; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2041 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_activate_5_T_4 ? buffer_3_47 : _GEN_2040; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2042 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_activate_5_T_4 ? buffer_3_48 : _GEN_2041; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2043 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_activate_5_T_4 ? buffer_3_49 : _GEN_2042; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2044 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_activate_5_T_4 ? buffer_3_50 : _GEN_2043; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2045 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_activate_5_T_4 ? buffer_3_51 : _GEN_2044; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2046 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_activate_5_T_4 ? buffer_3_52 : _GEN_2045; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2047 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_activate_5_T_4 ? buffer_3_53 : _GEN_2046; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2048 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_activate_5_T_4 ? buffer_3_54 : _GEN_2047; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2049 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_activate_5_T_4 ? buffer_3_55 : _GEN_2048; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2050 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_activate_5_T_4 ? buffer_3_56 : _GEN_2049; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2051 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_activate_5_T_4 ? buffer_3_57 : _GEN_2050; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2052 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_activate_5_T_4 ? buffer_3_58 : _GEN_2051; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2053 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_activate_5_T_4 ? buffer_3_59 : _GEN_2052; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2054 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_activate_5_T_4 ? buffer_3_60 : _GEN_2053; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2055 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_activate_5_T_4 ? buffer_3_61 : _GEN_2054; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2056 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_activate_5_T_4 ? buffer_3_62 : _GEN_2055; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2057 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_activate_5_T_4 ? buffer_3_63 : _GEN_2056; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2058 = 5'h5 < flow_ptr & flow_ptr <= 5'hd ? _GEN_2057 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [5:0] _io_out_activate_6_T_2 = 6'h30 + _io_out_activate_0_T_1; // @[Activation_Buffer.scala 76:88]
  wire [5:0] _io_out_activate_6_T_4 = _io_out_activate_6_T_2 - 6'h7; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_2060 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_activate_6_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2061 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_activate_6_T_4 ? buffer_0_2 : _GEN_2060; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2062 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_activate_6_T_4 ? buffer_0_3 : _GEN_2061; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2063 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_activate_6_T_4 ? buffer_0_4 : _GEN_2062; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2064 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_activate_6_T_4 ? buffer_0_5 : _GEN_2063; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2065 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_activate_6_T_4 ? buffer_0_6 : _GEN_2064; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2066 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_activate_6_T_4 ? buffer_0_7 : _GEN_2065; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2067 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_activate_6_T_4 ? buffer_0_8 : _GEN_2066; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2068 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_activate_6_T_4 ? buffer_0_9 : _GEN_2067; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2069 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_activate_6_T_4 ? buffer_0_10 : _GEN_2068; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2070 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_activate_6_T_4 ? buffer_0_11 : _GEN_2069; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2071 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_activate_6_T_4 ? buffer_0_12 : _GEN_2070; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2072 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_activate_6_T_4 ? buffer_0_13 : _GEN_2071; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2073 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_activate_6_T_4 ? buffer_0_14 : _GEN_2072; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2074 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_activate_6_T_4 ? buffer_0_15 : _GEN_2073; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2075 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_activate_6_T_4 ? buffer_0_16 : _GEN_2074; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2076 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_activate_6_T_4 ? buffer_0_17 : _GEN_2075; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2077 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_activate_6_T_4 ? buffer_0_18 : _GEN_2076; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2078 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_activate_6_T_4 ? buffer_0_19 : _GEN_2077; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2079 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_activate_6_T_4 ? buffer_0_20 : _GEN_2078; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2080 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_activate_6_T_4 ? buffer_0_21 : _GEN_2079; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2081 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_activate_6_T_4 ? buffer_0_22 : _GEN_2080; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2082 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_activate_6_T_4 ? buffer_0_23 : _GEN_2081; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2083 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_activate_6_T_4 ? buffer_0_24 : _GEN_2082; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2084 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_activate_6_T_4 ? buffer_0_25 : _GEN_2083; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2085 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_activate_6_T_4 ? buffer_0_26 : _GEN_2084; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2086 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_activate_6_T_4 ? buffer_0_27 : _GEN_2085; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2087 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_activate_6_T_4 ? buffer_0_28 : _GEN_2086; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2088 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_activate_6_T_4 ? buffer_0_29 : _GEN_2087; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2089 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_activate_6_T_4 ? buffer_0_30 : _GEN_2088; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2090 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_activate_6_T_4 ? buffer_0_31 : _GEN_2089; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2091 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_activate_6_T_4 ? buffer_0_32 : _GEN_2090; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2092 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_activate_6_T_4 ? buffer_0_33 : _GEN_2091; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2093 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_activate_6_T_4 ? buffer_0_34 : _GEN_2092; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2094 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_activate_6_T_4 ? buffer_0_35 : _GEN_2093; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2095 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_activate_6_T_4 ? buffer_0_36 : _GEN_2094; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2096 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_activate_6_T_4 ? buffer_0_37 : _GEN_2095; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2097 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_activate_6_T_4 ? buffer_0_38 : _GEN_2096; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2098 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_activate_6_T_4 ? buffer_0_39 : _GEN_2097; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2099 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_activate_6_T_4 ? buffer_0_40 : _GEN_2098; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2100 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_activate_6_T_4 ? buffer_0_41 : _GEN_2099; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2101 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_activate_6_T_4 ? buffer_0_42 : _GEN_2100; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2102 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_activate_6_T_4 ? buffer_0_43 : _GEN_2101; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2103 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_activate_6_T_4 ? buffer_0_44 : _GEN_2102; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2104 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_activate_6_T_4 ? buffer_0_45 : _GEN_2103; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2105 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_activate_6_T_4 ? buffer_0_46 : _GEN_2104; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2106 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_activate_6_T_4 ? buffer_0_47 : _GEN_2105; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2107 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_activate_6_T_4 ? buffer_0_48 : _GEN_2106; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2108 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_activate_6_T_4 ? buffer_0_49 : _GEN_2107; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2109 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_activate_6_T_4 ? buffer_0_50 : _GEN_2108; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2110 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_activate_6_T_4 ? buffer_0_51 : _GEN_2109; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2111 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_activate_6_T_4 ? buffer_0_52 : _GEN_2110; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2112 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_activate_6_T_4 ? buffer_0_53 : _GEN_2111; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2113 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_activate_6_T_4 ? buffer_0_54 : _GEN_2112; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2114 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_activate_6_T_4 ? buffer_0_55 : _GEN_2113; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2115 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_activate_6_T_4 ? buffer_0_56 : _GEN_2114; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2116 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_activate_6_T_4 ? buffer_0_57 : _GEN_2115; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2117 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_activate_6_T_4 ? buffer_0_58 : _GEN_2116; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2118 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_activate_6_T_4 ? buffer_0_59 : _GEN_2117; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2119 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_activate_6_T_4 ? buffer_0_60 : _GEN_2118; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2120 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_activate_6_T_4 ? buffer_0_61 : _GEN_2119; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2121 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_activate_6_T_4 ? buffer_0_62 : _GEN_2120; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2122 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_activate_6_T_4 ? buffer_0_63 : _GEN_2121; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2123 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_activate_6_T_4 ? buffer_1_0 : _GEN_2122; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2124 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_activate_6_T_4 ? buffer_1_1 : _GEN_2123; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2125 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_activate_6_T_4 ? buffer_1_2 : _GEN_2124; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2126 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_activate_6_T_4 ? buffer_1_3 : _GEN_2125; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2127 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_activate_6_T_4 ? buffer_1_4 : _GEN_2126; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2128 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_activate_6_T_4 ? buffer_1_5 : _GEN_2127; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2129 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_activate_6_T_4 ? buffer_1_6 : _GEN_2128; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2130 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_activate_6_T_4 ? buffer_1_7 : _GEN_2129; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2131 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_activate_6_T_4 ? buffer_1_8 : _GEN_2130; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2132 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_activate_6_T_4 ? buffer_1_9 : _GEN_2131; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2133 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_activate_6_T_4 ? buffer_1_10 : _GEN_2132; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2134 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_activate_6_T_4 ? buffer_1_11 : _GEN_2133; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2135 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_activate_6_T_4 ? buffer_1_12 : _GEN_2134; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2136 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_activate_6_T_4 ? buffer_1_13 : _GEN_2135; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2137 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_activate_6_T_4 ? buffer_1_14 : _GEN_2136; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2138 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_activate_6_T_4 ? buffer_1_15 : _GEN_2137; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2139 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_activate_6_T_4 ? buffer_1_16 : _GEN_2138; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2140 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_activate_6_T_4 ? buffer_1_17 : _GEN_2139; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2141 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_activate_6_T_4 ? buffer_1_18 : _GEN_2140; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2142 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_activate_6_T_4 ? buffer_1_19 : _GEN_2141; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2143 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_activate_6_T_4 ? buffer_1_20 : _GEN_2142; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2144 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_activate_6_T_4 ? buffer_1_21 : _GEN_2143; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2145 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_activate_6_T_4 ? buffer_1_22 : _GEN_2144; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2146 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_activate_6_T_4 ? buffer_1_23 : _GEN_2145; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2147 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_activate_6_T_4 ? buffer_1_24 : _GEN_2146; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2148 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_activate_6_T_4 ? buffer_1_25 : _GEN_2147; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2149 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_activate_6_T_4 ? buffer_1_26 : _GEN_2148; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2150 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_activate_6_T_4 ? buffer_1_27 : _GEN_2149; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2151 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_activate_6_T_4 ? buffer_1_28 : _GEN_2150; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2152 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_activate_6_T_4 ? buffer_1_29 : _GEN_2151; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2153 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_activate_6_T_4 ? buffer_1_30 : _GEN_2152; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2154 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_activate_6_T_4 ? buffer_1_31 : _GEN_2153; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2155 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_activate_6_T_4 ? buffer_1_32 : _GEN_2154; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2156 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_activate_6_T_4 ? buffer_1_33 : _GEN_2155; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2157 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_activate_6_T_4 ? buffer_1_34 : _GEN_2156; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2158 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_activate_6_T_4 ? buffer_1_35 : _GEN_2157; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2159 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_activate_6_T_4 ? buffer_1_36 : _GEN_2158; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2160 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_activate_6_T_4 ? buffer_1_37 : _GEN_2159; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2161 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_activate_6_T_4 ? buffer_1_38 : _GEN_2160; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2162 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_activate_6_T_4 ? buffer_1_39 : _GEN_2161; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2163 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_activate_6_T_4 ? buffer_1_40 : _GEN_2162; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2164 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_activate_6_T_4 ? buffer_1_41 : _GEN_2163; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2165 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_activate_6_T_4 ? buffer_1_42 : _GEN_2164; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2166 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_activate_6_T_4 ? buffer_1_43 : _GEN_2165; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2167 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_activate_6_T_4 ? buffer_1_44 : _GEN_2166; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2168 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_activate_6_T_4 ? buffer_1_45 : _GEN_2167; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2169 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_activate_6_T_4 ? buffer_1_46 : _GEN_2168; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2170 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_activate_6_T_4 ? buffer_1_47 : _GEN_2169; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2171 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_activate_6_T_4 ? buffer_1_48 : _GEN_2170; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2172 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_activate_6_T_4 ? buffer_1_49 : _GEN_2171; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2173 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_activate_6_T_4 ? buffer_1_50 : _GEN_2172; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2174 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_activate_6_T_4 ? buffer_1_51 : _GEN_2173; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2175 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_activate_6_T_4 ? buffer_1_52 : _GEN_2174; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2176 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_activate_6_T_4 ? buffer_1_53 : _GEN_2175; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2177 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_activate_6_T_4 ? buffer_1_54 : _GEN_2176; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2178 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_activate_6_T_4 ? buffer_1_55 : _GEN_2177; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2179 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_activate_6_T_4 ? buffer_1_56 : _GEN_2178; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2180 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_activate_6_T_4 ? buffer_1_57 : _GEN_2179; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2181 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_activate_6_T_4 ? buffer_1_58 : _GEN_2180; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2182 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_activate_6_T_4 ? buffer_1_59 : _GEN_2181; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2183 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_activate_6_T_4 ? buffer_1_60 : _GEN_2182; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2184 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_activate_6_T_4 ? buffer_1_61 : _GEN_2183; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2185 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_activate_6_T_4 ? buffer_1_62 : _GEN_2184; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2186 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_activate_6_T_4 ? buffer_1_63 : _GEN_2185; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2187 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_activate_6_T_4 ? buffer_2_0 : _GEN_2186; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2188 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_activate_6_T_4 ? buffer_2_1 : _GEN_2187; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2189 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_activate_6_T_4 ? buffer_2_2 : _GEN_2188; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2190 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_activate_6_T_4 ? buffer_2_3 : _GEN_2189; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2191 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_activate_6_T_4 ? buffer_2_4 : _GEN_2190; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2192 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_activate_6_T_4 ? buffer_2_5 : _GEN_2191; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2193 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_activate_6_T_4 ? buffer_2_6 : _GEN_2192; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2194 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_activate_6_T_4 ? buffer_2_7 : _GEN_2193; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2195 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_activate_6_T_4 ? buffer_2_8 : _GEN_2194; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2196 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_activate_6_T_4 ? buffer_2_9 : _GEN_2195; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2197 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_activate_6_T_4 ? buffer_2_10 : _GEN_2196; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2198 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_activate_6_T_4 ? buffer_2_11 : _GEN_2197; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2199 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_activate_6_T_4 ? buffer_2_12 : _GEN_2198; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2200 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_activate_6_T_4 ? buffer_2_13 : _GEN_2199; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2201 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_activate_6_T_4 ? buffer_2_14 : _GEN_2200; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2202 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_activate_6_T_4 ? buffer_2_15 : _GEN_2201; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2203 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_activate_6_T_4 ? buffer_2_16 : _GEN_2202; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2204 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_activate_6_T_4 ? buffer_2_17 : _GEN_2203; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2205 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_activate_6_T_4 ? buffer_2_18 : _GEN_2204; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2206 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_activate_6_T_4 ? buffer_2_19 : _GEN_2205; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2207 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_activate_6_T_4 ? buffer_2_20 : _GEN_2206; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2208 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_activate_6_T_4 ? buffer_2_21 : _GEN_2207; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2209 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_activate_6_T_4 ? buffer_2_22 : _GEN_2208; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2210 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_activate_6_T_4 ? buffer_2_23 : _GEN_2209; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2211 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_activate_6_T_4 ? buffer_2_24 : _GEN_2210; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2212 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_activate_6_T_4 ? buffer_2_25 : _GEN_2211; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2213 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_activate_6_T_4 ? buffer_2_26 : _GEN_2212; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2214 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_activate_6_T_4 ? buffer_2_27 : _GEN_2213; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2215 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_activate_6_T_4 ? buffer_2_28 : _GEN_2214; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2216 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_activate_6_T_4 ? buffer_2_29 : _GEN_2215; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2217 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_activate_6_T_4 ? buffer_2_30 : _GEN_2216; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2218 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_activate_6_T_4 ? buffer_2_31 : _GEN_2217; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2219 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_activate_6_T_4 ? buffer_2_32 : _GEN_2218; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2220 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_activate_6_T_4 ? buffer_2_33 : _GEN_2219; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2221 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_activate_6_T_4 ? buffer_2_34 : _GEN_2220; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2222 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_activate_6_T_4 ? buffer_2_35 : _GEN_2221; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2223 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_activate_6_T_4 ? buffer_2_36 : _GEN_2222; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2224 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_activate_6_T_4 ? buffer_2_37 : _GEN_2223; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2225 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_activate_6_T_4 ? buffer_2_38 : _GEN_2224; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2226 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_activate_6_T_4 ? buffer_2_39 : _GEN_2225; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2227 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_activate_6_T_4 ? buffer_2_40 : _GEN_2226; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2228 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_activate_6_T_4 ? buffer_2_41 : _GEN_2227; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2229 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_activate_6_T_4 ? buffer_2_42 : _GEN_2228; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2230 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_activate_6_T_4 ? buffer_2_43 : _GEN_2229; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2231 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_activate_6_T_4 ? buffer_2_44 : _GEN_2230; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2232 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_activate_6_T_4 ? buffer_2_45 : _GEN_2231; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2233 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_activate_6_T_4 ? buffer_2_46 : _GEN_2232; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2234 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_activate_6_T_4 ? buffer_2_47 : _GEN_2233; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2235 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_activate_6_T_4 ? buffer_2_48 : _GEN_2234; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2236 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_activate_6_T_4 ? buffer_2_49 : _GEN_2235; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2237 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_activate_6_T_4 ? buffer_2_50 : _GEN_2236; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2238 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_activate_6_T_4 ? buffer_2_51 : _GEN_2237; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2239 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_activate_6_T_4 ? buffer_2_52 : _GEN_2238; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2240 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_activate_6_T_4 ? buffer_2_53 : _GEN_2239; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2241 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_activate_6_T_4 ? buffer_2_54 : _GEN_2240; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2242 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_activate_6_T_4 ? buffer_2_55 : _GEN_2241; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2243 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_activate_6_T_4 ? buffer_2_56 : _GEN_2242; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2244 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_activate_6_T_4 ? buffer_2_57 : _GEN_2243; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2245 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_activate_6_T_4 ? buffer_2_58 : _GEN_2244; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2246 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_activate_6_T_4 ? buffer_2_59 : _GEN_2245; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2247 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_activate_6_T_4 ? buffer_2_60 : _GEN_2246; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2248 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_activate_6_T_4 ? buffer_2_61 : _GEN_2247; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2249 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_activate_6_T_4 ? buffer_2_62 : _GEN_2248; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2250 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_activate_6_T_4 ? buffer_2_63 : _GEN_2249; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2251 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_activate_6_T_4 ? buffer_3_0 : _GEN_2250; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2252 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_activate_6_T_4 ? buffer_3_1 : _GEN_2251; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2253 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_activate_6_T_4 ? buffer_3_2 : _GEN_2252; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2254 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_activate_6_T_4 ? buffer_3_3 : _GEN_2253; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2255 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_activate_6_T_4 ? buffer_3_4 : _GEN_2254; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2256 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_activate_6_T_4 ? buffer_3_5 : _GEN_2255; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2257 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_activate_6_T_4 ? buffer_3_6 : _GEN_2256; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2258 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_activate_6_T_4 ? buffer_3_7 : _GEN_2257; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2259 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_activate_6_T_4 ? buffer_3_8 : _GEN_2258; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2260 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_activate_6_T_4 ? buffer_3_9 : _GEN_2259; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2261 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_activate_6_T_4 ? buffer_3_10 : _GEN_2260; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2262 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_activate_6_T_4 ? buffer_3_11 : _GEN_2261; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2263 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_activate_6_T_4 ? buffer_3_12 : _GEN_2262; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2264 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_activate_6_T_4 ? buffer_3_13 : _GEN_2263; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2265 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_activate_6_T_4 ? buffer_3_14 : _GEN_2264; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2266 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_activate_6_T_4 ? buffer_3_15 : _GEN_2265; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2267 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_activate_6_T_4 ? buffer_3_16 : _GEN_2266; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2268 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_activate_6_T_4 ? buffer_3_17 : _GEN_2267; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2269 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_activate_6_T_4 ? buffer_3_18 : _GEN_2268; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2270 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_activate_6_T_4 ? buffer_3_19 : _GEN_2269; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2271 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_activate_6_T_4 ? buffer_3_20 : _GEN_2270; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2272 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_activate_6_T_4 ? buffer_3_21 : _GEN_2271; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2273 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_activate_6_T_4 ? buffer_3_22 : _GEN_2272; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2274 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_activate_6_T_4 ? buffer_3_23 : _GEN_2273; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2275 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_activate_6_T_4 ? buffer_3_24 : _GEN_2274; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2276 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_activate_6_T_4 ? buffer_3_25 : _GEN_2275; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2277 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_activate_6_T_4 ? buffer_3_26 : _GEN_2276; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2278 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_activate_6_T_4 ? buffer_3_27 : _GEN_2277; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2279 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_activate_6_T_4 ? buffer_3_28 : _GEN_2278; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2280 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_activate_6_T_4 ? buffer_3_29 : _GEN_2279; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2281 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_activate_6_T_4 ? buffer_3_30 : _GEN_2280; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2282 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_activate_6_T_4 ? buffer_3_31 : _GEN_2281; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2283 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_activate_6_T_4 ? buffer_3_32 : _GEN_2282; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2284 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_activate_6_T_4 ? buffer_3_33 : _GEN_2283; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2285 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_activate_6_T_4 ? buffer_3_34 : _GEN_2284; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2286 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_activate_6_T_4 ? buffer_3_35 : _GEN_2285; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2287 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_activate_6_T_4 ? buffer_3_36 : _GEN_2286; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2288 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_activate_6_T_4 ? buffer_3_37 : _GEN_2287; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2289 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_activate_6_T_4 ? buffer_3_38 : _GEN_2288; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2290 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_activate_6_T_4 ? buffer_3_39 : _GEN_2289; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2291 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_activate_6_T_4 ? buffer_3_40 : _GEN_2290; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2292 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_activate_6_T_4 ? buffer_3_41 : _GEN_2291; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2293 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_activate_6_T_4 ? buffer_3_42 : _GEN_2292; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2294 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_activate_6_T_4 ? buffer_3_43 : _GEN_2293; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2295 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_activate_6_T_4 ? buffer_3_44 : _GEN_2294; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2296 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_activate_6_T_4 ? buffer_3_45 : _GEN_2295; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2297 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_activate_6_T_4 ? buffer_3_46 : _GEN_2296; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2298 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_activate_6_T_4 ? buffer_3_47 : _GEN_2297; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2299 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_activate_6_T_4 ? buffer_3_48 : _GEN_2298; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2300 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_activate_6_T_4 ? buffer_3_49 : _GEN_2299; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2301 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_activate_6_T_4 ? buffer_3_50 : _GEN_2300; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2302 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_activate_6_T_4 ? buffer_3_51 : _GEN_2301; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2303 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_activate_6_T_4 ? buffer_3_52 : _GEN_2302; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2304 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_activate_6_T_4 ? buffer_3_53 : _GEN_2303; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2305 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_activate_6_T_4 ? buffer_3_54 : _GEN_2304; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2306 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_activate_6_T_4 ? buffer_3_55 : _GEN_2305; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2307 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_activate_6_T_4 ? buffer_3_56 : _GEN_2306; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2308 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_activate_6_T_4 ? buffer_3_57 : _GEN_2307; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2309 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_activate_6_T_4 ? buffer_3_58 : _GEN_2308; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2310 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_activate_6_T_4 ? buffer_3_59 : _GEN_2309; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2311 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_activate_6_T_4 ? buffer_3_60 : _GEN_2310; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2312 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_activate_6_T_4 ? buffer_3_61 : _GEN_2311; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2313 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_activate_6_T_4 ? buffer_3_62 : _GEN_2312; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2314 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_activate_6_T_4 ? buffer_3_63 : _GEN_2313; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2315 = 5'h6 < flow_ptr & flow_ptr <= 5'he ? _GEN_2314 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [5:0] _io_out_activate_7_T_2 = 6'h38 + _io_out_activate_0_T_1; // @[Activation_Buffer.scala 76:88]
  wire [5:0] _io_out_activate_7_T_4 = _io_out_activate_7_T_2 - 6'h8; // @[Activation_Buffer.scala 76:99]
  wire [7:0] _GEN_2317 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_activate_7_T_4 ? buffer_0_1 : buffer_0_0; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2318 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_activate_7_T_4 ? buffer_0_2 : _GEN_2317; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2319 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_activate_7_T_4 ? buffer_0_3 : _GEN_2318; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2320 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_activate_7_T_4 ? buffer_0_4 : _GEN_2319; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2321 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_activate_7_T_4 ? buffer_0_5 : _GEN_2320; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2322 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_activate_7_T_4 ? buffer_0_6 : _GEN_2321; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2323 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_activate_7_T_4 ? buffer_0_7 : _GEN_2322; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2324 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_activate_7_T_4 ? buffer_0_8 : _GEN_2323; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2325 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_activate_7_T_4 ? buffer_0_9 : _GEN_2324; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2326 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_activate_7_T_4 ? buffer_0_10 : _GEN_2325; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2327 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_activate_7_T_4 ? buffer_0_11 : _GEN_2326; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2328 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_activate_7_T_4 ? buffer_0_12 : _GEN_2327; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2329 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_activate_7_T_4 ? buffer_0_13 : _GEN_2328; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2330 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_activate_7_T_4 ? buffer_0_14 : _GEN_2329; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2331 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_activate_7_T_4 ? buffer_0_15 : _GEN_2330; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2332 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_activate_7_T_4 ? buffer_0_16 : _GEN_2331; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2333 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_activate_7_T_4 ? buffer_0_17 : _GEN_2332; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2334 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_activate_7_T_4 ? buffer_0_18 : _GEN_2333; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2335 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_activate_7_T_4 ? buffer_0_19 : _GEN_2334; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2336 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_activate_7_T_4 ? buffer_0_20 : _GEN_2335; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2337 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_activate_7_T_4 ? buffer_0_21 : _GEN_2336; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2338 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_activate_7_T_4 ? buffer_0_22 : _GEN_2337; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2339 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_activate_7_T_4 ? buffer_0_23 : _GEN_2338; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2340 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_activate_7_T_4 ? buffer_0_24 : _GEN_2339; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2341 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_activate_7_T_4 ? buffer_0_25 : _GEN_2340; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2342 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_activate_7_T_4 ? buffer_0_26 : _GEN_2341; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2343 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_activate_7_T_4 ? buffer_0_27 : _GEN_2342; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2344 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_activate_7_T_4 ? buffer_0_28 : _GEN_2343; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2345 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_activate_7_T_4 ? buffer_0_29 : _GEN_2344; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2346 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_activate_7_T_4 ? buffer_0_30 : _GEN_2345; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2347 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_activate_7_T_4 ? buffer_0_31 : _GEN_2346; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2348 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_activate_7_T_4 ? buffer_0_32 : _GEN_2347; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2349 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_activate_7_T_4 ? buffer_0_33 : _GEN_2348; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2350 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_activate_7_T_4 ? buffer_0_34 : _GEN_2349; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2351 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_activate_7_T_4 ? buffer_0_35 : _GEN_2350; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2352 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_activate_7_T_4 ? buffer_0_36 : _GEN_2351; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2353 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_activate_7_T_4 ? buffer_0_37 : _GEN_2352; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2354 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_activate_7_T_4 ? buffer_0_38 : _GEN_2353; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2355 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_activate_7_T_4 ? buffer_0_39 : _GEN_2354; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2356 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_activate_7_T_4 ? buffer_0_40 : _GEN_2355; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2357 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_activate_7_T_4 ? buffer_0_41 : _GEN_2356; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2358 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_activate_7_T_4 ? buffer_0_42 : _GEN_2357; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2359 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_activate_7_T_4 ? buffer_0_43 : _GEN_2358; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2360 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_activate_7_T_4 ? buffer_0_44 : _GEN_2359; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2361 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_activate_7_T_4 ? buffer_0_45 : _GEN_2360; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2362 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_activate_7_T_4 ? buffer_0_46 : _GEN_2361; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2363 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_activate_7_T_4 ? buffer_0_47 : _GEN_2362; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2364 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_activate_7_T_4 ? buffer_0_48 : _GEN_2363; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2365 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_activate_7_T_4 ? buffer_0_49 : _GEN_2364; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2366 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_activate_7_T_4 ? buffer_0_50 : _GEN_2365; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2367 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_activate_7_T_4 ? buffer_0_51 : _GEN_2366; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2368 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_activate_7_T_4 ? buffer_0_52 : _GEN_2367; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2369 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_activate_7_T_4 ? buffer_0_53 : _GEN_2368; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2370 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_activate_7_T_4 ? buffer_0_54 : _GEN_2369; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2371 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_activate_7_T_4 ? buffer_0_55 : _GEN_2370; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2372 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_activate_7_T_4 ? buffer_0_56 : _GEN_2371; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2373 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_activate_7_T_4 ? buffer_0_57 : _GEN_2372; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2374 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_activate_7_T_4 ? buffer_0_58 : _GEN_2373; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2375 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_activate_7_T_4 ? buffer_0_59 : _GEN_2374; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2376 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_activate_7_T_4 ? buffer_0_60 : _GEN_2375; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2377 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_activate_7_T_4 ? buffer_0_61 : _GEN_2376; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2378 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_activate_7_T_4 ? buffer_0_62 : _GEN_2377; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2379 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_activate_7_T_4 ? buffer_0_63 : _GEN_2378; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2380 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_activate_7_T_4 ? buffer_1_0 : _GEN_2379; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2381 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_activate_7_T_4 ? buffer_1_1 : _GEN_2380; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2382 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_activate_7_T_4 ? buffer_1_2 : _GEN_2381; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2383 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_activate_7_T_4 ? buffer_1_3 : _GEN_2382; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2384 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_activate_7_T_4 ? buffer_1_4 : _GEN_2383; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2385 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_activate_7_T_4 ? buffer_1_5 : _GEN_2384; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2386 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_activate_7_T_4 ? buffer_1_6 : _GEN_2385; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2387 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_activate_7_T_4 ? buffer_1_7 : _GEN_2386; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2388 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_activate_7_T_4 ? buffer_1_8 : _GEN_2387; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2389 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_activate_7_T_4 ? buffer_1_9 : _GEN_2388; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2390 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_activate_7_T_4 ? buffer_1_10 : _GEN_2389; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2391 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_activate_7_T_4 ? buffer_1_11 : _GEN_2390; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2392 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_activate_7_T_4 ? buffer_1_12 : _GEN_2391; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2393 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_activate_7_T_4 ? buffer_1_13 : _GEN_2392; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2394 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_activate_7_T_4 ? buffer_1_14 : _GEN_2393; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2395 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_activate_7_T_4 ? buffer_1_15 : _GEN_2394; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2396 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_activate_7_T_4 ? buffer_1_16 : _GEN_2395; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2397 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_activate_7_T_4 ? buffer_1_17 : _GEN_2396; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2398 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_activate_7_T_4 ? buffer_1_18 : _GEN_2397; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2399 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_activate_7_T_4 ? buffer_1_19 : _GEN_2398; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2400 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_activate_7_T_4 ? buffer_1_20 : _GEN_2399; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2401 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_activate_7_T_4 ? buffer_1_21 : _GEN_2400; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2402 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_activate_7_T_4 ? buffer_1_22 : _GEN_2401; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2403 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_activate_7_T_4 ? buffer_1_23 : _GEN_2402; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2404 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_activate_7_T_4 ? buffer_1_24 : _GEN_2403; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2405 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_activate_7_T_4 ? buffer_1_25 : _GEN_2404; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2406 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_activate_7_T_4 ? buffer_1_26 : _GEN_2405; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2407 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_activate_7_T_4 ? buffer_1_27 : _GEN_2406; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2408 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_activate_7_T_4 ? buffer_1_28 : _GEN_2407; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2409 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_activate_7_T_4 ? buffer_1_29 : _GEN_2408; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2410 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_activate_7_T_4 ? buffer_1_30 : _GEN_2409; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2411 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_activate_7_T_4 ? buffer_1_31 : _GEN_2410; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2412 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_activate_7_T_4 ? buffer_1_32 : _GEN_2411; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2413 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_activate_7_T_4 ? buffer_1_33 : _GEN_2412; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2414 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_activate_7_T_4 ? buffer_1_34 : _GEN_2413; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2415 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_activate_7_T_4 ? buffer_1_35 : _GEN_2414; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2416 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_activate_7_T_4 ? buffer_1_36 : _GEN_2415; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2417 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_activate_7_T_4 ? buffer_1_37 : _GEN_2416; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2418 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_activate_7_T_4 ? buffer_1_38 : _GEN_2417; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2419 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_activate_7_T_4 ? buffer_1_39 : _GEN_2418; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2420 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_activate_7_T_4 ? buffer_1_40 : _GEN_2419; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2421 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_activate_7_T_4 ? buffer_1_41 : _GEN_2420; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2422 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_activate_7_T_4 ? buffer_1_42 : _GEN_2421; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2423 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_activate_7_T_4 ? buffer_1_43 : _GEN_2422; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2424 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_activate_7_T_4 ? buffer_1_44 : _GEN_2423; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2425 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_activate_7_T_4 ? buffer_1_45 : _GEN_2424; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2426 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_activate_7_T_4 ? buffer_1_46 : _GEN_2425; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2427 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_activate_7_T_4 ? buffer_1_47 : _GEN_2426; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2428 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_activate_7_T_4 ? buffer_1_48 : _GEN_2427; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2429 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_activate_7_T_4 ? buffer_1_49 : _GEN_2428; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2430 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_activate_7_T_4 ? buffer_1_50 : _GEN_2429; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2431 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_activate_7_T_4 ? buffer_1_51 : _GEN_2430; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2432 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_activate_7_T_4 ? buffer_1_52 : _GEN_2431; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2433 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_activate_7_T_4 ? buffer_1_53 : _GEN_2432; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2434 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_activate_7_T_4 ? buffer_1_54 : _GEN_2433; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2435 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_activate_7_T_4 ? buffer_1_55 : _GEN_2434; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2436 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_activate_7_T_4 ? buffer_1_56 : _GEN_2435; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2437 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_activate_7_T_4 ? buffer_1_57 : _GEN_2436; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2438 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_activate_7_T_4 ? buffer_1_58 : _GEN_2437; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2439 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_activate_7_T_4 ? buffer_1_59 : _GEN_2438; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2440 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_activate_7_T_4 ? buffer_1_60 : _GEN_2439; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2441 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_activate_7_T_4 ? buffer_1_61 : _GEN_2440; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2442 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_activate_7_T_4 ? buffer_1_62 : _GEN_2441; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2443 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_activate_7_T_4 ? buffer_1_63 : _GEN_2442; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2444 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_activate_7_T_4 ? buffer_2_0 : _GEN_2443; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2445 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_activate_7_T_4 ? buffer_2_1 : _GEN_2444; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2446 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_activate_7_T_4 ? buffer_2_2 : _GEN_2445; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2447 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_activate_7_T_4 ? buffer_2_3 : _GEN_2446; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2448 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_activate_7_T_4 ? buffer_2_4 : _GEN_2447; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2449 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_activate_7_T_4 ? buffer_2_5 : _GEN_2448; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2450 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_activate_7_T_4 ? buffer_2_6 : _GEN_2449; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2451 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_activate_7_T_4 ? buffer_2_7 : _GEN_2450; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2452 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_activate_7_T_4 ? buffer_2_8 : _GEN_2451; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2453 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_activate_7_T_4 ? buffer_2_9 : _GEN_2452; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2454 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_activate_7_T_4 ? buffer_2_10 : _GEN_2453; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2455 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_activate_7_T_4 ? buffer_2_11 : _GEN_2454; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2456 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_activate_7_T_4 ? buffer_2_12 : _GEN_2455; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2457 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_activate_7_T_4 ? buffer_2_13 : _GEN_2456; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2458 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_activate_7_T_4 ? buffer_2_14 : _GEN_2457; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2459 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_activate_7_T_4 ? buffer_2_15 : _GEN_2458; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2460 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_activate_7_T_4 ? buffer_2_16 : _GEN_2459; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2461 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_activate_7_T_4 ? buffer_2_17 : _GEN_2460; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2462 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_activate_7_T_4 ? buffer_2_18 : _GEN_2461; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2463 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_activate_7_T_4 ? buffer_2_19 : _GEN_2462; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2464 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_activate_7_T_4 ? buffer_2_20 : _GEN_2463; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2465 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_activate_7_T_4 ? buffer_2_21 : _GEN_2464; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2466 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_activate_7_T_4 ? buffer_2_22 : _GEN_2465; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2467 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_activate_7_T_4 ? buffer_2_23 : _GEN_2466; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2468 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_activate_7_T_4 ? buffer_2_24 : _GEN_2467; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2469 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_activate_7_T_4 ? buffer_2_25 : _GEN_2468; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2470 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_activate_7_T_4 ? buffer_2_26 : _GEN_2469; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2471 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_activate_7_T_4 ? buffer_2_27 : _GEN_2470; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2472 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_activate_7_T_4 ? buffer_2_28 : _GEN_2471; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2473 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_activate_7_T_4 ? buffer_2_29 : _GEN_2472; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2474 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_activate_7_T_4 ? buffer_2_30 : _GEN_2473; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2475 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_activate_7_T_4 ? buffer_2_31 : _GEN_2474; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2476 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_activate_7_T_4 ? buffer_2_32 : _GEN_2475; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2477 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_activate_7_T_4 ? buffer_2_33 : _GEN_2476; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2478 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_activate_7_T_4 ? buffer_2_34 : _GEN_2477; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2479 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_activate_7_T_4 ? buffer_2_35 : _GEN_2478; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2480 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_activate_7_T_4 ? buffer_2_36 : _GEN_2479; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2481 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_activate_7_T_4 ? buffer_2_37 : _GEN_2480; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2482 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_activate_7_T_4 ? buffer_2_38 : _GEN_2481; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2483 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_activate_7_T_4 ? buffer_2_39 : _GEN_2482; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2484 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_activate_7_T_4 ? buffer_2_40 : _GEN_2483; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2485 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_activate_7_T_4 ? buffer_2_41 : _GEN_2484; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2486 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_activate_7_T_4 ? buffer_2_42 : _GEN_2485; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2487 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_activate_7_T_4 ? buffer_2_43 : _GEN_2486; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2488 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_activate_7_T_4 ? buffer_2_44 : _GEN_2487; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2489 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_activate_7_T_4 ? buffer_2_45 : _GEN_2488; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2490 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_activate_7_T_4 ? buffer_2_46 : _GEN_2489; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2491 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_activate_7_T_4 ? buffer_2_47 : _GEN_2490; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2492 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_activate_7_T_4 ? buffer_2_48 : _GEN_2491; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2493 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_activate_7_T_4 ? buffer_2_49 : _GEN_2492; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2494 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_activate_7_T_4 ? buffer_2_50 : _GEN_2493; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2495 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_activate_7_T_4 ? buffer_2_51 : _GEN_2494; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2496 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_activate_7_T_4 ? buffer_2_52 : _GEN_2495; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2497 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_activate_7_T_4 ? buffer_2_53 : _GEN_2496; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2498 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_activate_7_T_4 ? buffer_2_54 : _GEN_2497; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2499 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_activate_7_T_4 ? buffer_2_55 : _GEN_2498; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2500 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_activate_7_T_4 ? buffer_2_56 : _GEN_2499; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2501 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_activate_7_T_4 ? buffer_2_57 : _GEN_2500; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2502 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_activate_7_T_4 ? buffer_2_58 : _GEN_2501; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2503 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_activate_7_T_4 ? buffer_2_59 : _GEN_2502; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2504 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_activate_7_T_4 ? buffer_2_60 : _GEN_2503; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2505 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_activate_7_T_4 ? buffer_2_61 : _GEN_2504; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2506 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_activate_7_T_4 ? buffer_2_62 : _GEN_2505; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2507 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_activate_7_T_4 ? buffer_2_63 : _GEN_2506; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2508 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_activate_7_T_4 ? buffer_3_0 : _GEN_2507; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2509 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_activate_7_T_4 ? buffer_3_1 : _GEN_2508; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2510 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_activate_7_T_4 ? buffer_3_2 : _GEN_2509; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2511 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_activate_7_T_4 ? buffer_3_3 : _GEN_2510; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2512 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_activate_7_T_4 ? buffer_3_4 : _GEN_2511; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2513 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_activate_7_T_4 ? buffer_3_5 : _GEN_2512; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2514 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_activate_7_T_4 ? buffer_3_6 : _GEN_2513; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2515 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_activate_7_T_4 ? buffer_3_7 : _GEN_2514; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2516 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_activate_7_T_4 ? buffer_3_8 : _GEN_2515; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2517 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_activate_7_T_4 ? buffer_3_9 : _GEN_2516; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2518 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_activate_7_T_4 ? buffer_3_10 : _GEN_2517; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2519 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_activate_7_T_4 ? buffer_3_11 : _GEN_2518; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2520 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_activate_7_T_4 ? buffer_3_12 : _GEN_2519; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2521 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_activate_7_T_4 ? buffer_3_13 : _GEN_2520; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2522 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_activate_7_T_4 ? buffer_3_14 : _GEN_2521; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2523 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_activate_7_T_4 ? buffer_3_15 : _GEN_2522; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2524 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_activate_7_T_4 ? buffer_3_16 : _GEN_2523; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2525 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_activate_7_T_4 ? buffer_3_17 : _GEN_2524; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2526 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_activate_7_T_4 ? buffer_3_18 : _GEN_2525; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2527 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_activate_7_T_4 ? buffer_3_19 : _GEN_2526; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2528 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_activate_7_T_4 ? buffer_3_20 : _GEN_2527; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2529 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_activate_7_T_4 ? buffer_3_21 : _GEN_2528; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2530 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_activate_7_T_4 ? buffer_3_22 : _GEN_2529; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2531 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_activate_7_T_4 ? buffer_3_23 : _GEN_2530; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2532 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_activate_7_T_4 ? buffer_3_24 : _GEN_2531; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2533 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_activate_7_T_4 ? buffer_3_25 : _GEN_2532; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2534 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_activate_7_T_4 ? buffer_3_26 : _GEN_2533; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2535 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_activate_7_T_4 ? buffer_3_27 : _GEN_2534; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2536 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_activate_7_T_4 ? buffer_3_28 : _GEN_2535; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2537 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_activate_7_T_4 ? buffer_3_29 : _GEN_2536; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2538 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_activate_7_T_4 ? buffer_3_30 : _GEN_2537; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2539 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_activate_7_T_4 ? buffer_3_31 : _GEN_2538; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2540 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_activate_7_T_4 ? buffer_3_32 : _GEN_2539; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2541 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_activate_7_T_4 ? buffer_3_33 : _GEN_2540; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2542 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_activate_7_T_4 ? buffer_3_34 : _GEN_2541; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2543 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_activate_7_T_4 ? buffer_3_35 : _GEN_2542; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2544 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_activate_7_T_4 ? buffer_3_36 : _GEN_2543; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2545 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_activate_7_T_4 ? buffer_3_37 : _GEN_2544; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2546 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_activate_7_T_4 ? buffer_3_38 : _GEN_2545; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2547 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_activate_7_T_4 ? buffer_3_39 : _GEN_2546; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2548 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_activate_7_T_4 ? buffer_3_40 : _GEN_2547; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2549 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_activate_7_T_4 ? buffer_3_41 : _GEN_2548; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2550 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_activate_7_T_4 ? buffer_3_42 : _GEN_2549; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2551 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_activate_7_T_4 ? buffer_3_43 : _GEN_2550; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2552 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_activate_7_T_4 ? buffer_3_44 : _GEN_2551; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2553 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_activate_7_T_4 ? buffer_3_45 : _GEN_2552; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2554 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_activate_7_T_4 ? buffer_3_46 : _GEN_2553; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2555 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_activate_7_T_4 ? buffer_3_47 : _GEN_2554; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2556 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_activate_7_T_4 ? buffer_3_48 : _GEN_2555; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2557 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_activate_7_T_4 ? buffer_3_49 : _GEN_2556; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2558 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_activate_7_T_4 ? buffer_3_50 : _GEN_2557; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2559 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_activate_7_T_4 ? buffer_3_51 : _GEN_2558; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2560 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_activate_7_T_4 ? buffer_3_52 : _GEN_2559; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2561 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_activate_7_T_4 ? buffer_3_53 : _GEN_2560; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2562 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_activate_7_T_4 ? buffer_3_54 : _GEN_2561; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2563 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_activate_7_T_4 ? buffer_3_55 : _GEN_2562; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2564 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_activate_7_T_4 ? buffer_3_56 : _GEN_2563; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2565 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_activate_7_T_4 ? buffer_3_57 : _GEN_2564; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2566 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_activate_7_T_4 ? buffer_3_58 : _GEN_2565; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2567 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_activate_7_T_4 ? buffer_3_59 : _GEN_2566; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2568 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_activate_7_T_4 ? buffer_3_60 : _GEN_2567; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2569 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_activate_7_T_4 ? buffer_3_61 : _GEN_2568; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2570 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_activate_7_T_4 ? buffer_3_62 : _GEN_2569; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2571 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_activate_7_T_4 ? buffer_3_63 : _GEN_2570; // @[Activation_Buffer.scala 76:{28,28}]
  wire [7:0] _GEN_2572 = 5'h7 < flow_ptr & flow_ptr <= 5'hf ? _GEN_2571 : 8'h0; // @[Activation_Buffer.scala 75:65 76:28 78:28]
  wire [2:0] _read_ptr_T_1 = read_ptr + 3'h1; // @[Activation_Buffer.scala 88:26]
  assign io_out_activate_0 = _T_71 ? _GEN_773 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_1 = _T_71 ? _GEN_1030 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_2 = _T_71 ? _GEN_1287 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_3 = _T_71 ? _GEN_1544 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_4 = _T_71 ? _GEN_1801 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_5 = _T_71 ? _GEN_2058 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_6 = _T_71 ? _GEN_2315 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_activate_7 = _T_71 ? _GEN_2572 : 8'h0; // @[Activation_Buffer.scala 73:26 83:26]
  assign io_out_flow = flow_ptr != 5'h0; // @[Activation_Buffer.scala 67:17]
  assign io_isfull = read_ptr[1:0] == write_ptr[1:0] & read_ptr[2] != write_ptr[2]; // @[Activation_Buffer.scala 33:82]
  assign io_isempty = _full_T_2 & read_ptr[2] == write_ptr[2]; // @[Activation_Buffer.scala 34:83]
  assign io_isdone = flow_ptr == 5'h16; // @[Activation_Buffer.scala 93:17]
  always @(posedge clock) begin
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_0 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_0 <= io_in_data_x_0; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_1 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_1 <= io_in_data_x_8; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_2 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_2 <= io_in_data_x_16; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_3 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_3 <= io_in_data_x_24; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_4 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_4 <= io_in_data_x_32; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_5 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_5 <= io_in_data_x_40; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_6 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_6 <= io_in_data_x_48; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_7 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_7 <= io_in_data_x_56; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_8 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_8 <= io_in_data_x_1; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_9 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_9 <= io_in_data_x_9; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_10 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_10 <= io_in_data_x_17; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_11 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_11 <= io_in_data_x_25; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_12 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_12 <= io_in_data_x_33; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_13 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_13 <= io_in_data_x_41; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_14 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_14 <= io_in_data_x_49; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_15 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_15 <= io_in_data_x_57; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_16 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_16 <= io_in_data_x_2; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_17 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_17 <= io_in_data_x_10; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_18 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_18 <= io_in_data_x_18; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_19 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_19 <= io_in_data_x_26; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_20 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_20 <= io_in_data_x_34; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_21 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_21 <= io_in_data_x_42; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_22 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_22 <= io_in_data_x_50; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_23 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_23 <= io_in_data_x_58; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_24 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_24 <= io_in_data_x_3; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_25 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_25 <= io_in_data_x_11; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_26 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_26 <= io_in_data_x_19; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_27 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_27 <= io_in_data_x_27; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_28 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_28 <= io_in_data_x_35; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_29 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_29 <= io_in_data_x_43; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_30 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_30 <= io_in_data_x_51; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_31 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_31 <= io_in_data_x_59; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_32 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_32 <= io_in_data_x_4; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_33 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_33 <= io_in_data_x_12; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_34 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_34 <= io_in_data_x_20; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_35 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_35 <= io_in_data_x_28; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_36 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_36 <= io_in_data_x_36; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_37 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_37 <= io_in_data_x_44; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_38 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_38 <= io_in_data_x_52; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_39 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_39 <= io_in_data_x_60; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_40 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_40 <= io_in_data_x_5; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_41 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_41 <= io_in_data_x_13; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_42 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_42 <= io_in_data_x_21; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_43 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_43 <= io_in_data_x_29; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_44 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_44 <= io_in_data_x_37; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_45 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_45 <= io_in_data_x_45; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_46 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_46 <= io_in_data_x_53; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_47 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_47 <= io_in_data_x_61; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_48 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_48 <= io_in_data_x_6; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_49 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_49 <= io_in_data_x_14; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_50 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_50 <= io_in_data_x_22; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_51 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_51 <= io_in_data_x_30; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_52 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_52 <= io_in_data_x_38; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_53 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_53 <= io_in_data_x_46; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_54 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_54 <= io_in_data_x_54; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_55 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_55 <= io_in_data_x_62; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_56 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_56 <= io_in_data_x_7; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_57 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_57 <= io_in_data_x_15; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_58 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_58 <= io_in_data_x_23; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_59 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_59 <= io_in_data_x_31; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_60 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_60 <= io_in_data_x_39; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_61 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_61 <= io_in_data_x_47; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_62 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_62 <= io_in_data_x_55; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_0_63 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_0_63 <= io_in_data_x_63; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_0 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_0 <= io_in_data_x_0; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_1 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_1 <= io_in_data_x_8; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_2 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_2 <= io_in_data_x_16; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_3 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_3 <= io_in_data_x_24; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_4 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_4 <= io_in_data_x_32; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_5 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_5 <= io_in_data_x_40; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_6 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_6 <= io_in_data_x_48; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_7 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_7 <= io_in_data_x_56; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_8 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_8 <= io_in_data_x_1; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_9 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_9 <= io_in_data_x_9; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_10 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_10 <= io_in_data_x_17; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_11 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_11 <= io_in_data_x_25; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_12 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_12 <= io_in_data_x_33; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_13 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_13 <= io_in_data_x_41; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_14 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_14 <= io_in_data_x_49; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_15 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_15 <= io_in_data_x_57; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_16 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_16 <= io_in_data_x_2; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_17 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_17 <= io_in_data_x_10; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_18 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_18 <= io_in_data_x_18; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_19 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_19 <= io_in_data_x_26; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_20 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_20 <= io_in_data_x_34; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_21 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_21 <= io_in_data_x_42; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_22 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_22 <= io_in_data_x_50; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_23 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_23 <= io_in_data_x_58; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_24 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_24 <= io_in_data_x_3; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_25 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_25 <= io_in_data_x_11; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_26 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_26 <= io_in_data_x_19; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_27 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_27 <= io_in_data_x_27; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_28 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_28 <= io_in_data_x_35; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_29 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_29 <= io_in_data_x_43; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_30 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_30 <= io_in_data_x_51; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_31 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_31 <= io_in_data_x_59; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_32 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_32 <= io_in_data_x_4; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_33 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_33 <= io_in_data_x_12; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_34 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_34 <= io_in_data_x_20; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_35 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_35 <= io_in_data_x_28; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_36 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_36 <= io_in_data_x_36; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_37 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_37 <= io_in_data_x_44; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_38 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_38 <= io_in_data_x_52; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_39 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_39 <= io_in_data_x_60; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_40 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_40 <= io_in_data_x_5; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_41 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_41 <= io_in_data_x_13; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_42 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_42 <= io_in_data_x_21; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_43 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_43 <= io_in_data_x_29; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_44 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_44 <= io_in_data_x_37; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_45 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_45 <= io_in_data_x_45; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_46 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_46 <= io_in_data_x_53; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_47 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_47 <= io_in_data_x_61; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_48 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_48 <= io_in_data_x_6; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_49 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_49 <= io_in_data_x_14; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_50 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_50 <= io_in_data_x_22; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_51 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_51 <= io_in_data_x_30; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_52 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_52 <= io_in_data_x_38; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_53 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_53 <= io_in_data_x_46; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_54 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_54 <= io_in_data_x_54; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_55 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_55 <= io_in_data_x_62; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_56 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_56 <= io_in_data_x_7; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_57 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_57 <= io_in_data_x_15; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_58 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_58 <= io_in_data_x_23; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_59 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_59 <= io_in_data_x_31; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_60 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_60 <= io_in_data_x_39; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_61 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_61 <= io_in_data_x_47; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_62 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_62 <= io_in_data_x_55; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_1_63 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_1_63 <= io_in_data_x_63; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_0 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_0 <= io_in_data_x_0; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_1 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_1 <= io_in_data_x_8; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_2 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_2 <= io_in_data_x_16; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_3 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_3 <= io_in_data_x_24; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_4 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_4 <= io_in_data_x_32; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_5 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_5 <= io_in_data_x_40; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_6 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_6 <= io_in_data_x_48; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_7 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_7 <= io_in_data_x_56; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_8 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_8 <= io_in_data_x_1; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_9 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_9 <= io_in_data_x_9; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_10 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_10 <= io_in_data_x_17; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_11 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_11 <= io_in_data_x_25; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_12 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_12 <= io_in_data_x_33; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_13 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_13 <= io_in_data_x_41; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_14 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_14 <= io_in_data_x_49; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_15 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_15 <= io_in_data_x_57; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_16 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_16 <= io_in_data_x_2; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_17 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_17 <= io_in_data_x_10; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_18 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_18 <= io_in_data_x_18; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_19 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_19 <= io_in_data_x_26; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_20 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_20 <= io_in_data_x_34; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_21 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_21 <= io_in_data_x_42; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_22 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_22 <= io_in_data_x_50; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_23 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_23 <= io_in_data_x_58; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_24 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_24 <= io_in_data_x_3; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_25 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_25 <= io_in_data_x_11; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_26 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_26 <= io_in_data_x_19; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_27 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_27 <= io_in_data_x_27; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_28 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_28 <= io_in_data_x_35; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_29 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_29 <= io_in_data_x_43; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_30 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_30 <= io_in_data_x_51; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_31 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_31 <= io_in_data_x_59; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_32 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_32 <= io_in_data_x_4; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_33 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_33 <= io_in_data_x_12; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_34 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_34 <= io_in_data_x_20; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_35 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_35 <= io_in_data_x_28; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_36 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_36 <= io_in_data_x_36; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_37 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_37 <= io_in_data_x_44; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_38 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_38 <= io_in_data_x_52; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_39 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_39 <= io_in_data_x_60; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_40 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_40 <= io_in_data_x_5; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_41 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_41 <= io_in_data_x_13; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_42 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_42 <= io_in_data_x_21; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_43 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_43 <= io_in_data_x_29; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_44 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_44 <= io_in_data_x_37; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_45 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_45 <= io_in_data_x_45; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_46 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_46 <= io_in_data_x_53; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_47 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_47 <= io_in_data_x_61; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_48 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_48 <= io_in_data_x_6; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_49 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_49 <= io_in_data_x_14; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_50 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_50 <= io_in_data_x_22; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_51 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_51 <= io_in_data_x_30; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_52 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_52 <= io_in_data_x_38; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_53 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_53 <= io_in_data_x_46; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_54 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_54 <= io_in_data_x_54; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_55 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_55 <= io_in_data_x_62; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_56 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_56 <= io_in_data_x_7; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_57 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_57 <= io_in_data_x_15; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_58 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_58 <= io_in_data_x_23; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_59 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_59 <= io_in_data_x_31; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_60 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_60 <= io_in_data_x_39; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_61 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_61 <= io_in_data_x_47; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_62 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_62 <= io_in_data_x_55; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_2_63 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_2_63 <= io_in_data_x_63; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_0 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_0 <= io_in_data_x_0; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_1 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_1 <= io_in_data_x_8; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_2 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_2 <= io_in_data_x_16; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_3 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_3 <= io_in_data_x_24; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_4 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_4 <= io_in_data_x_32; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_5 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_5 <= io_in_data_x_40; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_6 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_6 <= io_in_data_x_48; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_7 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_7 <= io_in_data_x_56; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_8 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_8 <= io_in_data_x_1; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_9 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_9 <= io_in_data_x_9; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_10 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_10 <= io_in_data_x_17; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_11 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_11 <= io_in_data_x_25; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_12 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_12 <= io_in_data_x_33; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_13 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_13 <= io_in_data_x_41; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_14 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_14 <= io_in_data_x_49; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_15 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_15 <= io_in_data_x_57; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_16 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_16 <= io_in_data_x_2; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_17 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_17 <= io_in_data_x_10; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_18 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_18 <= io_in_data_x_18; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_19 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_19 <= io_in_data_x_26; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_20 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_20 <= io_in_data_x_34; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_21 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_21 <= io_in_data_x_42; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_22 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_22 <= io_in_data_x_50; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_23 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_23 <= io_in_data_x_58; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_24 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_24 <= io_in_data_x_3; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_25 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_25 <= io_in_data_x_11; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_26 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_26 <= io_in_data_x_19; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_27 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_27 <= io_in_data_x_27; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_28 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_28 <= io_in_data_x_35; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_29 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_29 <= io_in_data_x_43; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_30 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_30 <= io_in_data_x_51; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_31 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_31 <= io_in_data_x_59; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_32 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_32 <= io_in_data_x_4; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_33 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_33 <= io_in_data_x_12; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_34 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_34 <= io_in_data_x_20; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_35 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_35 <= io_in_data_x_28; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_36 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_36 <= io_in_data_x_36; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_37 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_37 <= io_in_data_x_44; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_38 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_38 <= io_in_data_x_52; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_39 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_39 <= io_in_data_x_60; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_40 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_40 <= io_in_data_x_5; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_41 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_41 <= io_in_data_x_13; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_42 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_42 <= io_in_data_x_21; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_43 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_43 <= io_in_data_x_29; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_44 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_44 <= io_in_data_x_37; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_45 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_45 <= io_in_data_x_45; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_46 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_46 <= io_in_data_x_53; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_47 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_47 <= io_in_data_x_61; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_48 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_48 <= io_in_data_x_6; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_49 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_49 <= io_in_data_x_14; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_50 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_50 <= io_in_data_x_22; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_51 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_51 <= io_in_data_x_30; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_52 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_52 <= io_in_data_x_38; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_53 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_53 <= io_in_data_x_46; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_54 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_54 <= io_in_data_x_54; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_55 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_55 <= io_in_data_x_62; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_56 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_56 <= io_in_data_x_7; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_57 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_57 <= io_in_data_x_15; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_58 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_58 <= io_in_data_x_23; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_59 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_59 <= io_in_data_x_31; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_60 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_60 <= io_in_data_x_39; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_61 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_61 <= io_in_data_x_47; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_62 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_62 <= io_in_data_x_55; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 24:23]
      buffer_3_63 <= 8'h0; // @[Activation_Buffer.scala 24:23]
    end else if (_T_1) begin // @[Activation_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Activation_Buffer.scala 49:68]
        buffer_3_63 <= io_in_data_x_63; // @[Activation_Buffer.scala 49:68]
      end
    end
    if (reset) begin // @[Activation_Buffer.scala 27:25]
      read_ptr <= 3'h0; // @[Activation_Buffer.scala 27:25]
    end else if (_T_70) begin // @[Activation_Buffer.scala 87:43]
      read_ptr <= _read_ptr_T_1; // @[Activation_Buffer.scala 88:14]
    end
    if (reset) begin // @[Activation_Buffer.scala 28:26]
      write_ptr <= 3'h0; // @[Activation_Buffer.scala 28:26]
    end else if (io_wen & ~full) begin // @[Activation_Buffer.scala 39:27]
      write_ptr <= _write_ptr_T_1; // @[Activation_Buffer.scala 40:15]
    end
    if (reset) begin // @[Activation_Buffer.scala 55:25]
      flow_ptr <= 5'h0; // @[Activation_Buffer.scala 55:25]
    end else if (io_ren & ~empty) begin // @[Activation_Buffer.scala 57:28]
      flow_ptr <= _flow_ptr_T_1; // @[Activation_Buffer.scala 58:14]
    end else if (flow_ptr == 5'h16) begin // @[Activation_Buffer.scala 59:49]
      flow_ptr <= 5'h0; // @[Activation_Buffer.scala 60:14]
    end else if (flow_ptr != 5'h0) begin // @[Activation_Buffer.scala 61:32]
      flow_ptr <= _flow_ptr_T_1; // @[Activation_Buffer.scala 62:14]
    end else begin
      flow_ptr <= 5'h0; // @[Activation_Buffer.scala 64:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buffer_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_0_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_0_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_0_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_0_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_0_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_0_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_0_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_0_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_0_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_0_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_0_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_0_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_0_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_0_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_0_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_0_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_0_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_0_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_0_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_0_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_0_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_0_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_0_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_0_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_0_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_0_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_0_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_0_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_0_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_0_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_0_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_0_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_0_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_0_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_0_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_0_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_0_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_0_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_0_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_0_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_0_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_0_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_0_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_0_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  buffer_0_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_0_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_0_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_0_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_0_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  buffer_0_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_0_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_0_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_0_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_0_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  buffer_0_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_0_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_0_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_0_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_0_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  buffer_1_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_1_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_1_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_1_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_1_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  buffer_1_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_1_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_1_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_1_8 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_1_9 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  buffer_1_10 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_1_11 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_1_12 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_1_13 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  buffer_1_14 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  buffer_1_15 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_1_16 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_1_17 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  buffer_1_18 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  buffer_1_19 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  buffer_1_20 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  buffer_1_21 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  buffer_1_22 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  buffer_1_23 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  buffer_1_24 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  buffer_1_25 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  buffer_1_26 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  buffer_1_27 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  buffer_1_28 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  buffer_1_29 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  buffer_1_30 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  buffer_1_31 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  buffer_1_32 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  buffer_1_33 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  buffer_1_34 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  buffer_1_35 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  buffer_1_36 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  buffer_1_37 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  buffer_1_38 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  buffer_1_39 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  buffer_1_40 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  buffer_1_41 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  buffer_1_42 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  buffer_1_43 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  buffer_1_44 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  buffer_1_45 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  buffer_1_46 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  buffer_1_47 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  buffer_1_48 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  buffer_1_49 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  buffer_1_50 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  buffer_1_51 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  buffer_1_52 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  buffer_1_53 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  buffer_1_54 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  buffer_1_55 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  buffer_1_56 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  buffer_1_57 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  buffer_1_58 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  buffer_1_59 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  buffer_1_60 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  buffer_1_61 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  buffer_1_62 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  buffer_1_63 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  buffer_2_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  buffer_2_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  buffer_2_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  buffer_2_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  buffer_2_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  buffer_2_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  buffer_2_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  buffer_2_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  buffer_2_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  buffer_2_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  buffer_2_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  buffer_2_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  buffer_2_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  buffer_2_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  buffer_2_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  buffer_2_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  buffer_2_16 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  buffer_2_17 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  buffer_2_18 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  buffer_2_19 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  buffer_2_20 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  buffer_2_21 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  buffer_2_22 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  buffer_2_23 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  buffer_2_24 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  buffer_2_25 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  buffer_2_26 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  buffer_2_27 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  buffer_2_28 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  buffer_2_29 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  buffer_2_30 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  buffer_2_31 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  buffer_2_32 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  buffer_2_33 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  buffer_2_34 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  buffer_2_35 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  buffer_2_36 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  buffer_2_37 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  buffer_2_38 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  buffer_2_39 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  buffer_2_40 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  buffer_2_41 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  buffer_2_42 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  buffer_2_43 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  buffer_2_44 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  buffer_2_45 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  buffer_2_46 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  buffer_2_47 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  buffer_2_48 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  buffer_2_49 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  buffer_2_50 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  buffer_2_51 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  buffer_2_52 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  buffer_2_53 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  buffer_2_54 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  buffer_2_55 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  buffer_2_56 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  buffer_2_57 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  buffer_2_58 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  buffer_2_59 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  buffer_2_60 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  buffer_2_61 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  buffer_2_62 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  buffer_2_63 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  buffer_3_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  buffer_3_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  buffer_3_2 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  buffer_3_3 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  buffer_3_4 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  buffer_3_5 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  buffer_3_6 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  buffer_3_7 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  buffer_3_8 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  buffer_3_9 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  buffer_3_10 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  buffer_3_11 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  buffer_3_12 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  buffer_3_13 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  buffer_3_14 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  buffer_3_15 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  buffer_3_16 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  buffer_3_17 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  buffer_3_18 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  buffer_3_19 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  buffer_3_20 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  buffer_3_21 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  buffer_3_22 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  buffer_3_23 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  buffer_3_24 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  buffer_3_25 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  buffer_3_26 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  buffer_3_27 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  buffer_3_28 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  buffer_3_29 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  buffer_3_30 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  buffer_3_31 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  buffer_3_32 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  buffer_3_33 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  buffer_3_34 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  buffer_3_35 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  buffer_3_36 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  buffer_3_37 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  buffer_3_38 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  buffer_3_39 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  buffer_3_40 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  buffer_3_41 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  buffer_3_42 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  buffer_3_43 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  buffer_3_44 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  buffer_3_45 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  buffer_3_46 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  buffer_3_47 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  buffer_3_48 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  buffer_3_49 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  buffer_3_50 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  buffer_3_51 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  buffer_3_52 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  buffer_3_53 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  buffer_3_54 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  buffer_3_55 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  buffer_3_56 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  buffer_3_57 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  buffer_3_58 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  buffer_3_59 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  buffer_3_60 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  buffer_3_61 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  buffer_3_62 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  buffer_3_63 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  read_ptr = _RAND_256[2:0];
  _RAND_257 = {1{`RANDOM}};
  write_ptr = _RAND_257[2:0];
  _RAND_258 = {1{`RANDOM}};
  flow_ptr = _RAND_258[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Weight_Buffer(
  input        clock,
  input        reset,
  input        io_wen,
  input        io_ren,
  input  [7:0] io_in_weight_x_0,
  input  [7:0] io_in_weight_x_1,
  input  [7:0] io_in_weight_x_2,
  input  [7:0] io_in_weight_x_3,
  input  [7:0] io_in_weight_x_4,
  input  [7:0] io_in_weight_x_5,
  input  [7:0] io_in_weight_x_6,
  input  [7:0] io_in_weight_x_7,
  input  [7:0] io_in_weight_x_8,
  input  [7:0] io_in_weight_x_9,
  input  [7:0] io_in_weight_x_10,
  input  [7:0] io_in_weight_x_11,
  input  [7:0] io_in_weight_x_12,
  input  [7:0] io_in_weight_x_13,
  input  [7:0] io_in_weight_x_14,
  input  [7:0] io_in_weight_x_15,
  input  [7:0] io_in_weight_x_16,
  input  [7:0] io_in_weight_x_17,
  input  [7:0] io_in_weight_x_18,
  input  [7:0] io_in_weight_x_19,
  input  [7:0] io_in_weight_x_20,
  input  [7:0] io_in_weight_x_21,
  input  [7:0] io_in_weight_x_22,
  input  [7:0] io_in_weight_x_23,
  input  [7:0] io_in_weight_x_24,
  input  [7:0] io_in_weight_x_25,
  input  [7:0] io_in_weight_x_26,
  input  [7:0] io_in_weight_x_27,
  input  [7:0] io_in_weight_x_28,
  input  [7:0] io_in_weight_x_29,
  input  [7:0] io_in_weight_x_30,
  input  [7:0] io_in_weight_x_31,
  input  [7:0] io_in_weight_x_32,
  input  [7:0] io_in_weight_x_33,
  input  [7:0] io_in_weight_x_34,
  input  [7:0] io_in_weight_x_35,
  input  [7:0] io_in_weight_x_36,
  input  [7:0] io_in_weight_x_37,
  input  [7:0] io_in_weight_x_38,
  input  [7:0] io_in_weight_x_39,
  input  [7:0] io_in_weight_x_40,
  input  [7:0] io_in_weight_x_41,
  input  [7:0] io_in_weight_x_42,
  input  [7:0] io_in_weight_x_43,
  input  [7:0] io_in_weight_x_44,
  input  [7:0] io_in_weight_x_45,
  input  [7:0] io_in_weight_x_46,
  input  [7:0] io_in_weight_x_47,
  input  [7:0] io_in_weight_x_48,
  input  [7:0] io_in_weight_x_49,
  input  [7:0] io_in_weight_x_50,
  input  [7:0] io_in_weight_x_51,
  input  [7:0] io_in_weight_x_52,
  input  [7:0] io_in_weight_x_53,
  input  [7:0] io_in_weight_x_54,
  input  [7:0] io_in_weight_x_55,
  input  [7:0] io_in_weight_x_56,
  input  [7:0] io_in_weight_x_57,
  input  [7:0] io_in_weight_x_58,
  input  [7:0] io_in_weight_x_59,
  input  [7:0] io_in_weight_x_60,
  input  [7:0] io_in_weight_x_61,
  input  [7:0] io_in_weight_x_62,
  input  [7:0] io_in_weight_x_63,
  output [7:0] io_out_weight_0,
  output [7:0] io_out_weight_1,
  output [7:0] io_out_weight_2,
  output [7:0] io_out_weight_3,
  output [7:0] io_out_weight_4,
  output [7:0] io_out_weight_5,
  output [7:0] io_out_weight_6,
  output [7:0] io_out_weight_7,
  output       io_out_shift,
  output       io_isfull,
  output       io_isempty,
  output       io_isdone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] buffer_0_0; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_1; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_2; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_3; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_4; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_5; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_6; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_7; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_8; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_9; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_10; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_11; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_12; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_13; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_14; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_15; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_16; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_17; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_18; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_19; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_20; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_21; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_22; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_23; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_24; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_25; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_26; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_27; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_28; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_29; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_30; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_31; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_32; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_33; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_34; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_35; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_36; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_37; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_38; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_39; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_40; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_41; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_42; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_43; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_44; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_45; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_46; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_47; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_48; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_49; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_50; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_51; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_52; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_53; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_54; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_55; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_56; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_57; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_58; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_59; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_60; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_61; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_62; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_0_63; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_0; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_1; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_2; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_3; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_4; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_5; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_6; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_7; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_8; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_9; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_10; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_11; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_12; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_13; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_14; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_15; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_16; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_17; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_18; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_19; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_20; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_21; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_22; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_23; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_24; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_25; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_26; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_27; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_28; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_29; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_30; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_31; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_32; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_33; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_34; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_35; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_36; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_37; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_38; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_39; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_40; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_41; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_42; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_43; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_44; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_45; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_46; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_47; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_48; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_49; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_50; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_51; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_52; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_53; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_54; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_55; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_56; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_57; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_58; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_59; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_60; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_61; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_62; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_1_63; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_0; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_1; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_2; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_3; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_4; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_5; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_6; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_7; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_8; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_9; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_10; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_11; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_12; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_13; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_14; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_15; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_16; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_17; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_18; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_19; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_20; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_21; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_22; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_23; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_24; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_25; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_26; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_27; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_28; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_29; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_30; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_31; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_32; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_33; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_34; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_35; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_36; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_37; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_38; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_39; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_40; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_41; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_42; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_43; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_44; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_45; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_46; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_47; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_48; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_49; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_50; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_51; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_52; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_53; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_54; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_55; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_56; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_57; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_58; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_59; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_60; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_61; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_62; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_2_63; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_0; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_1; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_2; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_3; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_4; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_5; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_6; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_7; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_8; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_9; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_10; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_11; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_12; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_13; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_14; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_15; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_16; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_17; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_18; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_19; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_20; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_21; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_22; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_23; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_24; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_25; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_26; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_27; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_28; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_29; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_30; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_31; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_32; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_33; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_34; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_35; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_36; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_37; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_38; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_39; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_40; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_41; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_42; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_43; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_44; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_45; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_46; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_47; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_48; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_49; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_50; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_51; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_52; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_53; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_54; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_55; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_56; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_57; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_58; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_59; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_60; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_61; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_62; // @[Weight_Buffer.scala 25:23]
  reg [7:0] buffer_3_63; // @[Weight_Buffer.scala 25:23]
  reg [2:0] read_ptr; // @[Weight_Buffer.scala 28:25]
  reg [2:0] write_ptr; // @[Weight_Buffer.scala 29:26]
  wire  _full_T_2 = read_ptr[1:0] == write_ptr[1:0]; // @[Weight_Buffer.scala 34:42]
  wire  full = read_ptr[1:0] == write_ptr[1:0] & read_ptr[2] != write_ptr[2]; // @[Weight_Buffer.scala 34:78]
  wire  empty = _full_T_2 & read_ptr[2] == write_ptr[2]; // @[Weight_Buffer.scala 35:79]
  wire  _T_1 = io_wen & ~full; // @[Weight_Buffer.scala 40:15]
  wire [2:0] _write_ptr_T_1 = write_ptr + 3'h1; // @[Weight_Buffer.scala 41:28]
  reg [3:0] shift_ptr; // @[Weight_Buffer.scala 51:26]
  wire [3:0] _shift_ptr_T_1 = shift_ptr - 4'h1; // @[Weight_Buffer.scala 54:28]
  wire [7:0] _io_out_weight_0_T_1 = shift_ptr * 4'h8; // @[Weight_Buffer.scala 64:75]
  wire [8:0] _io_out_weight_0_T_2 = {{1'd0}, _io_out_weight_0_T_1}; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_516 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_0_T_2[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_517 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_0_T_2[5:0] ? buffer_0_2 : _GEN_516; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_518 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_0_T_2[5:0] ? buffer_0_3 : _GEN_517; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_519 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_0_T_2[5:0] ? buffer_0_4 : _GEN_518; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_520 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_0_T_2[5:0] ? buffer_0_5 : _GEN_519; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_521 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_0_T_2[5:0] ? buffer_0_6 : _GEN_520; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_522 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_0_T_2[5:0] ? buffer_0_7 : _GEN_521; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_523 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_0_T_2[5:0] ? buffer_0_8 : _GEN_522; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_524 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_0_T_2[5:0] ? buffer_0_9 : _GEN_523; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_525 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_0_T_2[5:0] ? buffer_0_10 : _GEN_524; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_526 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_0_T_2[5:0] ? buffer_0_11 : _GEN_525; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_527 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_0_T_2[5:0] ? buffer_0_12 : _GEN_526; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_528 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_0_T_2[5:0] ? buffer_0_13 : _GEN_527; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_529 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_0_T_2[5:0] ? buffer_0_14 : _GEN_528; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_530 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_0_T_2[5:0] ? buffer_0_15 : _GEN_529; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_531 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_0_T_2[5:0] ? buffer_0_16 : _GEN_530; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_532 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_0_T_2[5:0] ? buffer_0_17 : _GEN_531; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_533 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_0_T_2[5:0] ? buffer_0_18 : _GEN_532; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_534 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_0_T_2[5:0] ? buffer_0_19 : _GEN_533; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_535 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_0_T_2[5:0] ? buffer_0_20 : _GEN_534; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_536 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_0_T_2[5:0] ? buffer_0_21 : _GEN_535; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_537 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_0_T_2[5:0] ? buffer_0_22 : _GEN_536; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_538 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_0_T_2[5:0] ? buffer_0_23 : _GEN_537; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_539 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_0_T_2[5:0] ? buffer_0_24 : _GEN_538; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_540 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_0_T_2[5:0] ? buffer_0_25 : _GEN_539; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_541 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_0_T_2[5:0] ? buffer_0_26 : _GEN_540; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_542 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_0_T_2[5:0] ? buffer_0_27 : _GEN_541; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_543 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_0_T_2[5:0] ? buffer_0_28 : _GEN_542; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_544 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_0_T_2[5:0] ? buffer_0_29 : _GEN_543; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_545 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_0_T_2[5:0] ? buffer_0_30 : _GEN_544; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_546 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_0_T_2[5:0] ? buffer_0_31 : _GEN_545; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_547 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_0_T_2[5:0] ? buffer_0_32 : _GEN_546; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_548 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_0_T_2[5:0] ? buffer_0_33 : _GEN_547; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_549 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_0_T_2[5:0] ? buffer_0_34 : _GEN_548; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_550 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_0_T_2[5:0] ? buffer_0_35 : _GEN_549; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_551 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_0_T_2[5:0] ? buffer_0_36 : _GEN_550; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_552 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_0_T_2[5:0] ? buffer_0_37 : _GEN_551; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_553 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_0_T_2[5:0] ? buffer_0_38 : _GEN_552; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_554 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_0_T_2[5:0] ? buffer_0_39 : _GEN_553; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_555 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_0_T_2[5:0] ? buffer_0_40 : _GEN_554; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_556 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_0_T_2[5:0] ? buffer_0_41 : _GEN_555; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_557 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_0_T_2[5:0] ? buffer_0_42 : _GEN_556; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_558 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_0_T_2[5:0] ? buffer_0_43 : _GEN_557; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_559 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_0_T_2[5:0] ? buffer_0_44 : _GEN_558; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_560 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_0_T_2[5:0] ? buffer_0_45 : _GEN_559; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_561 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_0_T_2[5:0] ? buffer_0_46 : _GEN_560; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_562 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_0_T_2[5:0] ? buffer_0_47 : _GEN_561; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_563 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_0_T_2[5:0] ? buffer_0_48 : _GEN_562; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_564 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_0_T_2[5:0] ? buffer_0_49 : _GEN_563; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_565 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_0_T_2[5:0] ? buffer_0_50 : _GEN_564; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_566 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_0_T_2[5:0] ? buffer_0_51 : _GEN_565; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_567 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_0_T_2[5:0] ? buffer_0_52 : _GEN_566; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_568 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_0_T_2[5:0] ? buffer_0_53 : _GEN_567; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_569 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_0_T_2[5:0] ? buffer_0_54 : _GEN_568; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_570 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_0_T_2[5:0] ? buffer_0_55 : _GEN_569; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_571 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_0_T_2[5:0] ? buffer_0_56 : _GEN_570; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_572 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_0_T_2[5:0] ? buffer_0_57 : _GEN_571; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_573 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_0_T_2[5:0] ? buffer_0_58 : _GEN_572; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_574 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_0_T_2[5:0] ? buffer_0_59 : _GEN_573; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_575 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_0_T_2[5:0] ? buffer_0_60 : _GEN_574; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_576 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_0_T_2[5:0] ? buffer_0_61 : _GEN_575; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_577 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_0_T_2[5:0] ? buffer_0_62 : _GEN_576; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_578 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_0_T_2[5:0] ? buffer_0_63 : _GEN_577; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_579 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_0_T_2[5:0] ? buffer_1_0 : _GEN_578; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_580 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_0_T_2[5:0] ? buffer_1_1 : _GEN_579; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_581 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_0_T_2[5:0] ? buffer_1_2 : _GEN_580; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_582 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_0_T_2[5:0] ? buffer_1_3 : _GEN_581; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_583 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_0_T_2[5:0] ? buffer_1_4 : _GEN_582; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_584 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_0_T_2[5:0] ? buffer_1_5 : _GEN_583; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_585 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_0_T_2[5:0] ? buffer_1_6 : _GEN_584; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_586 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_0_T_2[5:0] ? buffer_1_7 : _GEN_585; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_587 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_0_T_2[5:0] ? buffer_1_8 : _GEN_586; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_588 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_0_T_2[5:0] ? buffer_1_9 : _GEN_587; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_589 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_0_T_2[5:0] ? buffer_1_10 : _GEN_588; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_590 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_0_T_2[5:0] ? buffer_1_11 : _GEN_589; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_591 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_0_T_2[5:0] ? buffer_1_12 : _GEN_590; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_592 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_0_T_2[5:0] ? buffer_1_13 : _GEN_591; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_593 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_0_T_2[5:0] ? buffer_1_14 : _GEN_592; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_594 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_0_T_2[5:0] ? buffer_1_15 : _GEN_593; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_595 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_0_T_2[5:0] ? buffer_1_16 : _GEN_594; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_596 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_0_T_2[5:0] ? buffer_1_17 : _GEN_595; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_597 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_0_T_2[5:0] ? buffer_1_18 : _GEN_596; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_598 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_0_T_2[5:0] ? buffer_1_19 : _GEN_597; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_599 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_0_T_2[5:0] ? buffer_1_20 : _GEN_598; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_600 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_0_T_2[5:0] ? buffer_1_21 : _GEN_599; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_601 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_0_T_2[5:0] ? buffer_1_22 : _GEN_600; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_602 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_0_T_2[5:0] ? buffer_1_23 : _GEN_601; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_603 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_0_T_2[5:0] ? buffer_1_24 : _GEN_602; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_604 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_0_T_2[5:0] ? buffer_1_25 : _GEN_603; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_605 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_0_T_2[5:0] ? buffer_1_26 : _GEN_604; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_606 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_0_T_2[5:0] ? buffer_1_27 : _GEN_605; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_607 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_0_T_2[5:0] ? buffer_1_28 : _GEN_606; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_608 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_0_T_2[5:0] ? buffer_1_29 : _GEN_607; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_609 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_0_T_2[5:0] ? buffer_1_30 : _GEN_608; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_610 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_0_T_2[5:0] ? buffer_1_31 : _GEN_609; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_611 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_0_T_2[5:0] ? buffer_1_32 : _GEN_610; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_612 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_0_T_2[5:0] ? buffer_1_33 : _GEN_611; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_613 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_0_T_2[5:0] ? buffer_1_34 : _GEN_612; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_614 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_0_T_2[5:0] ? buffer_1_35 : _GEN_613; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_615 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_0_T_2[5:0] ? buffer_1_36 : _GEN_614; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_616 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_0_T_2[5:0] ? buffer_1_37 : _GEN_615; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_617 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_0_T_2[5:0] ? buffer_1_38 : _GEN_616; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_618 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_0_T_2[5:0] ? buffer_1_39 : _GEN_617; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_619 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_0_T_2[5:0] ? buffer_1_40 : _GEN_618; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_620 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_0_T_2[5:0] ? buffer_1_41 : _GEN_619; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_621 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_0_T_2[5:0] ? buffer_1_42 : _GEN_620; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_622 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_0_T_2[5:0] ? buffer_1_43 : _GEN_621; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_623 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_0_T_2[5:0] ? buffer_1_44 : _GEN_622; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_624 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_0_T_2[5:0] ? buffer_1_45 : _GEN_623; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_625 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_0_T_2[5:0] ? buffer_1_46 : _GEN_624; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_626 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_0_T_2[5:0] ? buffer_1_47 : _GEN_625; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_627 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_0_T_2[5:0] ? buffer_1_48 : _GEN_626; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_628 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_0_T_2[5:0] ? buffer_1_49 : _GEN_627; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_629 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_0_T_2[5:0] ? buffer_1_50 : _GEN_628; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_630 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_0_T_2[5:0] ? buffer_1_51 : _GEN_629; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_631 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_0_T_2[5:0] ? buffer_1_52 : _GEN_630; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_632 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_0_T_2[5:0] ? buffer_1_53 : _GEN_631; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_633 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_0_T_2[5:0] ? buffer_1_54 : _GEN_632; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_634 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_0_T_2[5:0] ? buffer_1_55 : _GEN_633; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_635 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_0_T_2[5:0] ? buffer_1_56 : _GEN_634; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_636 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_0_T_2[5:0] ? buffer_1_57 : _GEN_635; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_637 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_0_T_2[5:0] ? buffer_1_58 : _GEN_636; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_638 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_0_T_2[5:0] ? buffer_1_59 : _GEN_637; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_639 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_0_T_2[5:0] ? buffer_1_60 : _GEN_638; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_640 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_0_T_2[5:0] ? buffer_1_61 : _GEN_639; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_641 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_0_T_2[5:0] ? buffer_1_62 : _GEN_640; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_642 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_0_T_2[5:0] ? buffer_1_63 : _GEN_641; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_643 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_0_T_2[5:0] ? buffer_2_0 : _GEN_642; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_644 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_0_T_2[5:0] ? buffer_2_1 : _GEN_643; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_645 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_0_T_2[5:0] ? buffer_2_2 : _GEN_644; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_646 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_0_T_2[5:0] ? buffer_2_3 : _GEN_645; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_647 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_0_T_2[5:0] ? buffer_2_4 : _GEN_646; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_648 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_0_T_2[5:0] ? buffer_2_5 : _GEN_647; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_649 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_0_T_2[5:0] ? buffer_2_6 : _GEN_648; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_650 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_0_T_2[5:0] ? buffer_2_7 : _GEN_649; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_651 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_0_T_2[5:0] ? buffer_2_8 : _GEN_650; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_652 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_0_T_2[5:0] ? buffer_2_9 : _GEN_651; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_653 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_0_T_2[5:0] ? buffer_2_10 : _GEN_652; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_654 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_0_T_2[5:0] ? buffer_2_11 : _GEN_653; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_655 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_0_T_2[5:0] ? buffer_2_12 : _GEN_654; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_656 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_0_T_2[5:0] ? buffer_2_13 : _GEN_655; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_657 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_0_T_2[5:0] ? buffer_2_14 : _GEN_656; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_658 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_0_T_2[5:0] ? buffer_2_15 : _GEN_657; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_659 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_0_T_2[5:0] ? buffer_2_16 : _GEN_658; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_660 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_0_T_2[5:0] ? buffer_2_17 : _GEN_659; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_661 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_0_T_2[5:0] ? buffer_2_18 : _GEN_660; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_662 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_0_T_2[5:0] ? buffer_2_19 : _GEN_661; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_663 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_0_T_2[5:0] ? buffer_2_20 : _GEN_662; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_664 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_0_T_2[5:0] ? buffer_2_21 : _GEN_663; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_665 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_0_T_2[5:0] ? buffer_2_22 : _GEN_664; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_666 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_0_T_2[5:0] ? buffer_2_23 : _GEN_665; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_667 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_0_T_2[5:0] ? buffer_2_24 : _GEN_666; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_668 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_0_T_2[5:0] ? buffer_2_25 : _GEN_667; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_669 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_0_T_2[5:0] ? buffer_2_26 : _GEN_668; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_670 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_0_T_2[5:0] ? buffer_2_27 : _GEN_669; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_671 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_0_T_2[5:0] ? buffer_2_28 : _GEN_670; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_672 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_0_T_2[5:0] ? buffer_2_29 : _GEN_671; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_673 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_0_T_2[5:0] ? buffer_2_30 : _GEN_672; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_674 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_0_T_2[5:0] ? buffer_2_31 : _GEN_673; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_675 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_0_T_2[5:0] ? buffer_2_32 : _GEN_674; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_676 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_0_T_2[5:0] ? buffer_2_33 : _GEN_675; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_677 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_0_T_2[5:0] ? buffer_2_34 : _GEN_676; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_678 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_0_T_2[5:0] ? buffer_2_35 : _GEN_677; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_679 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_0_T_2[5:0] ? buffer_2_36 : _GEN_678; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_680 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_0_T_2[5:0] ? buffer_2_37 : _GEN_679; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_681 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_0_T_2[5:0] ? buffer_2_38 : _GEN_680; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_682 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_0_T_2[5:0] ? buffer_2_39 : _GEN_681; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_683 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_0_T_2[5:0] ? buffer_2_40 : _GEN_682; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_684 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_0_T_2[5:0] ? buffer_2_41 : _GEN_683; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_685 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_0_T_2[5:0] ? buffer_2_42 : _GEN_684; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_686 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_0_T_2[5:0] ? buffer_2_43 : _GEN_685; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_687 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_0_T_2[5:0] ? buffer_2_44 : _GEN_686; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_688 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_0_T_2[5:0] ? buffer_2_45 : _GEN_687; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_689 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_0_T_2[5:0] ? buffer_2_46 : _GEN_688; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_690 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_0_T_2[5:0] ? buffer_2_47 : _GEN_689; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_691 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_0_T_2[5:0] ? buffer_2_48 : _GEN_690; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_692 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_0_T_2[5:0] ? buffer_2_49 : _GEN_691; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_693 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_0_T_2[5:0] ? buffer_2_50 : _GEN_692; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_694 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_0_T_2[5:0] ? buffer_2_51 : _GEN_693; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_695 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_0_T_2[5:0] ? buffer_2_52 : _GEN_694; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_696 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_0_T_2[5:0] ? buffer_2_53 : _GEN_695; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_697 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_0_T_2[5:0] ? buffer_2_54 : _GEN_696; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_698 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_0_T_2[5:0] ? buffer_2_55 : _GEN_697; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_699 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_0_T_2[5:0] ? buffer_2_56 : _GEN_698; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_700 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_0_T_2[5:0] ? buffer_2_57 : _GEN_699; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_701 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_0_T_2[5:0] ? buffer_2_58 : _GEN_700; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_702 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_0_T_2[5:0] ? buffer_2_59 : _GEN_701; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_703 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_0_T_2[5:0] ? buffer_2_60 : _GEN_702; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_704 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_0_T_2[5:0] ? buffer_2_61 : _GEN_703; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_705 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_0_T_2[5:0] ? buffer_2_62 : _GEN_704; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_706 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_0_T_2[5:0] ? buffer_2_63 : _GEN_705; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_707 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_0_T_2[5:0] ? buffer_3_0 : _GEN_706; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_708 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_0_T_2[5:0] ? buffer_3_1 : _GEN_707; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_709 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_0_T_2[5:0] ? buffer_3_2 : _GEN_708; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_710 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_0_T_2[5:0] ? buffer_3_3 : _GEN_709; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_711 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_0_T_2[5:0] ? buffer_3_4 : _GEN_710; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_712 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_0_T_2[5:0] ? buffer_3_5 : _GEN_711; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_713 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_0_T_2[5:0] ? buffer_3_6 : _GEN_712; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_714 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_0_T_2[5:0] ? buffer_3_7 : _GEN_713; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_715 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_0_T_2[5:0] ? buffer_3_8 : _GEN_714; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_716 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_0_T_2[5:0] ? buffer_3_9 : _GEN_715; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_717 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_0_T_2[5:0] ? buffer_3_10 : _GEN_716; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_718 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_0_T_2[5:0] ? buffer_3_11 : _GEN_717; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_719 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_0_T_2[5:0] ? buffer_3_12 : _GEN_718; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_720 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_0_T_2[5:0] ? buffer_3_13 : _GEN_719; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_721 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_0_T_2[5:0] ? buffer_3_14 : _GEN_720; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_722 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_0_T_2[5:0] ? buffer_3_15 : _GEN_721; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_723 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_0_T_2[5:0] ? buffer_3_16 : _GEN_722; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_724 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_0_T_2[5:0] ? buffer_3_17 : _GEN_723; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_725 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_0_T_2[5:0] ? buffer_3_18 : _GEN_724; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_726 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_0_T_2[5:0] ? buffer_3_19 : _GEN_725; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_727 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_0_T_2[5:0] ? buffer_3_20 : _GEN_726; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_728 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_0_T_2[5:0] ? buffer_3_21 : _GEN_727; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_729 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_0_T_2[5:0] ? buffer_3_22 : _GEN_728; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_730 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_0_T_2[5:0] ? buffer_3_23 : _GEN_729; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_731 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_0_T_2[5:0] ? buffer_3_24 : _GEN_730; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_732 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_0_T_2[5:0] ? buffer_3_25 : _GEN_731; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_733 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_0_T_2[5:0] ? buffer_3_26 : _GEN_732; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_734 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_0_T_2[5:0] ? buffer_3_27 : _GEN_733; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_735 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_0_T_2[5:0] ? buffer_3_28 : _GEN_734; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_736 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_0_T_2[5:0] ? buffer_3_29 : _GEN_735; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_737 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_0_T_2[5:0] ? buffer_3_30 : _GEN_736; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_738 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_0_T_2[5:0] ? buffer_3_31 : _GEN_737; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_739 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_0_T_2[5:0] ? buffer_3_32 : _GEN_738; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_740 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_0_T_2[5:0] ? buffer_3_33 : _GEN_739; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_741 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_0_T_2[5:0] ? buffer_3_34 : _GEN_740; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_742 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_0_T_2[5:0] ? buffer_3_35 : _GEN_741; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_743 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_0_T_2[5:0] ? buffer_3_36 : _GEN_742; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_744 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_0_T_2[5:0] ? buffer_3_37 : _GEN_743; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_745 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_0_T_2[5:0] ? buffer_3_38 : _GEN_744; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_746 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_0_T_2[5:0] ? buffer_3_39 : _GEN_745; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_747 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_0_T_2[5:0] ? buffer_3_40 : _GEN_746; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_748 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_0_T_2[5:0] ? buffer_3_41 : _GEN_747; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_749 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_0_T_2[5:0] ? buffer_3_42 : _GEN_748; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_750 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_0_T_2[5:0] ? buffer_3_43 : _GEN_749; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_751 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_0_T_2[5:0] ? buffer_3_44 : _GEN_750; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_752 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_0_T_2[5:0] ? buffer_3_45 : _GEN_751; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_753 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_0_T_2[5:0] ? buffer_3_46 : _GEN_752; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_754 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_0_T_2[5:0] ? buffer_3_47 : _GEN_753; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_755 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_0_T_2[5:0] ? buffer_3_48 : _GEN_754; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_756 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_0_T_2[5:0] ? buffer_3_49 : _GEN_755; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_757 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_0_T_2[5:0] ? buffer_3_50 : _GEN_756; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_758 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_0_T_2[5:0] ? buffer_3_51 : _GEN_757; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_759 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_0_T_2[5:0] ? buffer_3_52 : _GEN_758; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_760 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_0_T_2[5:0] ? buffer_3_53 : _GEN_759; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_761 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_0_T_2[5:0] ? buffer_3_54 : _GEN_760; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_762 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_0_T_2[5:0] ? buffer_3_55 : _GEN_761; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_763 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_0_T_2[5:0] ? buffer_3_56 : _GEN_762; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_764 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_0_T_2[5:0] ? buffer_3_57 : _GEN_763; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_765 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_0_T_2[5:0] ? buffer_3_58 : _GEN_764; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_766 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_0_T_2[5:0] ? buffer_3_59 : _GEN_765; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_767 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_0_T_2[5:0] ? buffer_3_60 : _GEN_766; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_768 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_0_T_2[5:0] ? buffer_3_61 : _GEN_767; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_769 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_0_T_2[5:0] ? buffer_3_62 : _GEN_768; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_770 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_0_T_2[5:0] ? buffer_3_63 : _GEN_769; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_1_T_3 = _io_out_weight_0_T_1 + 8'h1; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_772 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_1_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_773 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_1_T_3[5:0] ? buffer_0_2 : _GEN_772; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_774 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_1_T_3[5:0] ? buffer_0_3 : _GEN_773; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_775 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_1_T_3[5:0] ? buffer_0_4 : _GEN_774; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_776 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_1_T_3[5:0] ? buffer_0_5 : _GEN_775; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_777 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_1_T_3[5:0] ? buffer_0_6 : _GEN_776; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_778 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_1_T_3[5:0] ? buffer_0_7 : _GEN_777; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_779 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_1_T_3[5:0] ? buffer_0_8 : _GEN_778; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_780 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_1_T_3[5:0] ? buffer_0_9 : _GEN_779; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_781 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_1_T_3[5:0] ? buffer_0_10 : _GEN_780; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_782 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_1_T_3[5:0] ? buffer_0_11 : _GEN_781; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_783 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_1_T_3[5:0] ? buffer_0_12 : _GEN_782; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_784 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_1_T_3[5:0] ? buffer_0_13 : _GEN_783; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_785 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_1_T_3[5:0] ? buffer_0_14 : _GEN_784; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_786 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_1_T_3[5:0] ? buffer_0_15 : _GEN_785; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_787 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_1_T_3[5:0] ? buffer_0_16 : _GEN_786; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_788 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_1_T_3[5:0] ? buffer_0_17 : _GEN_787; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_789 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_1_T_3[5:0] ? buffer_0_18 : _GEN_788; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_790 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_1_T_3[5:0] ? buffer_0_19 : _GEN_789; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_791 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_1_T_3[5:0] ? buffer_0_20 : _GEN_790; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_792 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_1_T_3[5:0] ? buffer_0_21 : _GEN_791; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_793 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_1_T_3[5:0] ? buffer_0_22 : _GEN_792; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_794 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_1_T_3[5:0] ? buffer_0_23 : _GEN_793; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_795 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_1_T_3[5:0] ? buffer_0_24 : _GEN_794; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_796 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_1_T_3[5:0] ? buffer_0_25 : _GEN_795; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_797 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_1_T_3[5:0] ? buffer_0_26 : _GEN_796; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_798 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_1_T_3[5:0] ? buffer_0_27 : _GEN_797; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_799 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_1_T_3[5:0] ? buffer_0_28 : _GEN_798; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_800 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_1_T_3[5:0] ? buffer_0_29 : _GEN_799; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_801 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_1_T_3[5:0] ? buffer_0_30 : _GEN_800; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_802 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_1_T_3[5:0] ? buffer_0_31 : _GEN_801; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_803 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_1_T_3[5:0] ? buffer_0_32 : _GEN_802; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_804 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_1_T_3[5:0] ? buffer_0_33 : _GEN_803; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_805 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_1_T_3[5:0] ? buffer_0_34 : _GEN_804; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_806 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_1_T_3[5:0] ? buffer_0_35 : _GEN_805; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_807 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_1_T_3[5:0] ? buffer_0_36 : _GEN_806; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_808 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_1_T_3[5:0] ? buffer_0_37 : _GEN_807; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_809 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_1_T_3[5:0] ? buffer_0_38 : _GEN_808; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_810 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_1_T_3[5:0] ? buffer_0_39 : _GEN_809; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_811 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_1_T_3[5:0] ? buffer_0_40 : _GEN_810; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_812 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_1_T_3[5:0] ? buffer_0_41 : _GEN_811; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_813 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_1_T_3[5:0] ? buffer_0_42 : _GEN_812; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_814 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_1_T_3[5:0] ? buffer_0_43 : _GEN_813; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_815 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_1_T_3[5:0] ? buffer_0_44 : _GEN_814; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_816 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_1_T_3[5:0] ? buffer_0_45 : _GEN_815; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_817 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_1_T_3[5:0] ? buffer_0_46 : _GEN_816; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_818 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_1_T_3[5:0] ? buffer_0_47 : _GEN_817; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_819 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_1_T_3[5:0] ? buffer_0_48 : _GEN_818; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_820 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_1_T_3[5:0] ? buffer_0_49 : _GEN_819; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_821 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_1_T_3[5:0] ? buffer_0_50 : _GEN_820; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_822 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_1_T_3[5:0] ? buffer_0_51 : _GEN_821; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_823 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_1_T_3[5:0] ? buffer_0_52 : _GEN_822; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_824 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_1_T_3[5:0] ? buffer_0_53 : _GEN_823; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_825 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_1_T_3[5:0] ? buffer_0_54 : _GEN_824; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_826 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_1_T_3[5:0] ? buffer_0_55 : _GEN_825; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_827 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_1_T_3[5:0] ? buffer_0_56 : _GEN_826; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_828 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_1_T_3[5:0] ? buffer_0_57 : _GEN_827; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_829 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_1_T_3[5:0] ? buffer_0_58 : _GEN_828; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_830 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_1_T_3[5:0] ? buffer_0_59 : _GEN_829; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_831 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_1_T_3[5:0] ? buffer_0_60 : _GEN_830; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_832 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_1_T_3[5:0] ? buffer_0_61 : _GEN_831; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_833 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_1_T_3[5:0] ? buffer_0_62 : _GEN_832; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_834 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_1_T_3[5:0] ? buffer_0_63 : _GEN_833; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_835 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_1_T_3[5:0] ? buffer_1_0 : _GEN_834; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_836 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_1_T_3[5:0] ? buffer_1_1 : _GEN_835; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_837 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_1_T_3[5:0] ? buffer_1_2 : _GEN_836; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_838 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_1_T_3[5:0] ? buffer_1_3 : _GEN_837; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_839 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_1_T_3[5:0] ? buffer_1_4 : _GEN_838; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_840 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_1_T_3[5:0] ? buffer_1_5 : _GEN_839; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_841 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_1_T_3[5:0] ? buffer_1_6 : _GEN_840; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_842 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_1_T_3[5:0] ? buffer_1_7 : _GEN_841; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_843 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_1_T_3[5:0] ? buffer_1_8 : _GEN_842; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_844 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_1_T_3[5:0] ? buffer_1_9 : _GEN_843; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_845 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_1_T_3[5:0] ? buffer_1_10 : _GEN_844; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_846 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_1_T_3[5:0] ? buffer_1_11 : _GEN_845; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_847 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_1_T_3[5:0] ? buffer_1_12 : _GEN_846; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_848 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_1_T_3[5:0] ? buffer_1_13 : _GEN_847; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_849 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_1_T_3[5:0] ? buffer_1_14 : _GEN_848; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_850 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_1_T_3[5:0] ? buffer_1_15 : _GEN_849; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_851 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_1_T_3[5:0] ? buffer_1_16 : _GEN_850; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_852 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_1_T_3[5:0] ? buffer_1_17 : _GEN_851; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_853 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_1_T_3[5:0] ? buffer_1_18 : _GEN_852; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_854 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_1_T_3[5:0] ? buffer_1_19 : _GEN_853; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_855 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_1_T_3[5:0] ? buffer_1_20 : _GEN_854; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_856 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_1_T_3[5:0] ? buffer_1_21 : _GEN_855; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_857 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_1_T_3[5:0] ? buffer_1_22 : _GEN_856; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_858 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_1_T_3[5:0] ? buffer_1_23 : _GEN_857; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_859 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_1_T_3[5:0] ? buffer_1_24 : _GEN_858; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_860 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_1_T_3[5:0] ? buffer_1_25 : _GEN_859; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_861 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_1_T_3[5:0] ? buffer_1_26 : _GEN_860; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_862 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_1_T_3[5:0] ? buffer_1_27 : _GEN_861; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_863 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_1_T_3[5:0] ? buffer_1_28 : _GEN_862; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_864 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_1_T_3[5:0] ? buffer_1_29 : _GEN_863; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_865 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_1_T_3[5:0] ? buffer_1_30 : _GEN_864; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_866 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_1_T_3[5:0] ? buffer_1_31 : _GEN_865; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_867 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_1_T_3[5:0] ? buffer_1_32 : _GEN_866; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_868 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_1_T_3[5:0] ? buffer_1_33 : _GEN_867; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_869 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_1_T_3[5:0] ? buffer_1_34 : _GEN_868; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_870 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_1_T_3[5:0] ? buffer_1_35 : _GEN_869; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_871 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_1_T_3[5:0] ? buffer_1_36 : _GEN_870; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_872 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_1_T_3[5:0] ? buffer_1_37 : _GEN_871; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_873 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_1_T_3[5:0] ? buffer_1_38 : _GEN_872; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_874 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_1_T_3[5:0] ? buffer_1_39 : _GEN_873; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_875 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_1_T_3[5:0] ? buffer_1_40 : _GEN_874; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_876 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_1_T_3[5:0] ? buffer_1_41 : _GEN_875; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_877 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_1_T_3[5:0] ? buffer_1_42 : _GEN_876; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_878 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_1_T_3[5:0] ? buffer_1_43 : _GEN_877; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_879 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_1_T_3[5:0] ? buffer_1_44 : _GEN_878; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_880 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_1_T_3[5:0] ? buffer_1_45 : _GEN_879; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_881 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_1_T_3[5:0] ? buffer_1_46 : _GEN_880; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_882 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_1_T_3[5:0] ? buffer_1_47 : _GEN_881; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_883 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_1_T_3[5:0] ? buffer_1_48 : _GEN_882; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_884 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_1_T_3[5:0] ? buffer_1_49 : _GEN_883; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_885 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_1_T_3[5:0] ? buffer_1_50 : _GEN_884; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_886 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_1_T_3[5:0] ? buffer_1_51 : _GEN_885; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_887 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_1_T_3[5:0] ? buffer_1_52 : _GEN_886; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_888 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_1_T_3[5:0] ? buffer_1_53 : _GEN_887; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_889 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_1_T_3[5:0] ? buffer_1_54 : _GEN_888; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_890 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_1_T_3[5:0] ? buffer_1_55 : _GEN_889; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_891 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_1_T_3[5:0] ? buffer_1_56 : _GEN_890; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_892 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_1_T_3[5:0] ? buffer_1_57 : _GEN_891; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_893 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_1_T_3[5:0] ? buffer_1_58 : _GEN_892; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_894 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_1_T_3[5:0] ? buffer_1_59 : _GEN_893; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_895 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_1_T_3[5:0] ? buffer_1_60 : _GEN_894; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_896 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_1_T_3[5:0] ? buffer_1_61 : _GEN_895; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_897 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_1_T_3[5:0] ? buffer_1_62 : _GEN_896; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_898 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_1_T_3[5:0] ? buffer_1_63 : _GEN_897; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_899 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_1_T_3[5:0] ? buffer_2_0 : _GEN_898; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_900 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_1_T_3[5:0] ? buffer_2_1 : _GEN_899; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_901 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_1_T_3[5:0] ? buffer_2_2 : _GEN_900; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_902 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_1_T_3[5:0] ? buffer_2_3 : _GEN_901; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_903 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_1_T_3[5:0] ? buffer_2_4 : _GEN_902; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_904 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_1_T_3[5:0] ? buffer_2_5 : _GEN_903; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_905 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_1_T_3[5:0] ? buffer_2_6 : _GEN_904; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_906 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_1_T_3[5:0] ? buffer_2_7 : _GEN_905; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_907 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_1_T_3[5:0] ? buffer_2_8 : _GEN_906; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_908 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_1_T_3[5:0] ? buffer_2_9 : _GEN_907; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_909 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_1_T_3[5:0] ? buffer_2_10 : _GEN_908; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_910 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_1_T_3[5:0] ? buffer_2_11 : _GEN_909; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_911 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_1_T_3[5:0] ? buffer_2_12 : _GEN_910; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_912 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_1_T_3[5:0] ? buffer_2_13 : _GEN_911; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_913 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_1_T_3[5:0] ? buffer_2_14 : _GEN_912; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_914 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_1_T_3[5:0] ? buffer_2_15 : _GEN_913; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_915 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_1_T_3[5:0] ? buffer_2_16 : _GEN_914; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_916 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_1_T_3[5:0] ? buffer_2_17 : _GEN_915; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_917 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_1_T_3[5:0] ? buffer_2_18 : _GEN_916; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_918 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_1_T_3[5:0] ? buffer_2_19 : _GEN_917; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_919 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_1_T_3[5:0] ? buffer_2_20 : _GEN_918; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_920 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_1_T_3[5:0] ? buffer_2_21 : _GEN_919; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_921 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_1_T_3[5:0] ? buffer_2_22 : _GEN_920; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_922 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_1_T_3[5:0] ? buffer_2_23 : _GEN_921; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_923 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_1_T_3[5:0] ? buffer_2_24 : _GEN_922; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_924 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_1_T_3[5:0] ? buffer_2_25 : _GEN_923; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_925 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_1_T_3[5:0] ? buffer_2_26 : _GEN_924; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_926 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_1_T_3[5:0] ? buffer_2_27 : _GEN_925; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_927 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_1_T_3[5:0] ? buffer_2_28 : _GEN_926; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_928 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_1_T_3[5:0] ? buffer_2_29 : _GEN_927; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_929 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_1_T_3[5:0] ? buffer_2_30 : _GEN_928; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_930 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_1_T_3[5:0] ? buffer_2_31 : _GEN_929; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_931 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_1_T_3[5:0] ? buffer_2_32 : _GEN_930; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_932 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_1_T_3[5:0] ? buffer_2_33 : _GEN_931; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_933 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_1_T_3[5:0] ? buffer_2_34 : _GEN_932; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_934 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_1_T_3[5:0] ? buffer_2_35 : _GEN_933; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_935 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_1_T_3[5:0] ? buffer_2_36 : _GEN_934; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_936 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_1_T_3[5:0] ? buffer_2_37 : _GEN_935; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_937 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_1_T_3[5:0] ? buffer_2_38 : _GEN_936; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_938 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_1_T_3[5:0] ? buffer_2_39 : _GEN_937; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_939 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_1_T_3[5:0] ? buffer_2_40 : _GEN_938; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_940 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_1_T_3[5:0] ? buffer_2_41 : _GEN_939; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_941 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_1_T_3[5:0] ? buffer_2_42 : _GEN_940; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_942 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_1_T_3[5:0] ? buffer_2_43 : _GEN_941; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_943 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_1_T_3[5:0] ? buffer_2_44 : _GEN_942; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_944 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_1_T_3[5:0] ? buffer_2_45 : _GEN_943; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_945 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_1_T_3[5:0] ? buffer_2_46 : _GEN_944; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_946 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_1_T_3[5:0] ? buffer_2_47 : _GEN_945; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_947 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_1_T_3[5:0] ? buffer_2_48 : _GEN_946; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_948 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_1_T_3[5:0] ? buffer_2_49 : _GEN_947; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_949 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_1_T_3[5:0] ? buffer_2_50 : _GEN_948; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_950 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_1_T_3[5:0] ? buffer_2_51 : _GEN_949; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_951 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_1_T_3[5:0] ? buffer_2_52 : _GEN_950; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_952 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_1_T_3[5:0] ? buffer_2_53 : _GEN_951; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_953 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_1_T_3[5:0] ? buffer_2_54 : _GEN_952; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_954 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_1_T_3[5:0] ? buffer_2_55 : _GEN_953; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_955 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_1_T_3[5:0] ? buffer_2_56 : _GEN_954; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_956 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_1_T_3[5:0] ? buffer_2_57 : _GEN_955; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_957 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_1_T_3[5:0] ? buffer_2_58 : _GEN_956; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_958 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_1_T_3[5:0] ? buffer_2_59 : _GEN_957; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_959 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_1_T_3[5:0] ? buffer_2_60 : _GEN_958; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_960 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_1_T_3[5:0] ? buffer_2_61 : _GEN_959; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_961 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_1_T_3[5:0] ? buffer_2_62 : _GEN_960; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_962 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_1_T_3[5:0] ? buffer_2_63 : _GEN_961; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_963 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_1_T_3[5:0] ? buffer_3_0 : _GEN_962; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_964 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_1_T_3[5:0] ? buffer_3_1 : _GEN_963; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_965 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_1_T_3[5:0] ? buffer_3_2 : _GEN_964; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_966 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_1_T_3[5:0] ? buffer_3_3 : _GEN_965; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_967 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_1_T_3[5:0] ? buffer_3_4 : _GEN_966; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_968 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_1_T_3[5:0] ? buffer_3_5 : _GEN_967; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_969 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_1_T_3[5:0] ? buffer_3_6 : _GEN_968; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_970 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_1_T_3[5:0] ? buffer_3_7 : _GEN_969; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_971 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_1_T_3[5:0] ? buffer_3_8 : _GEN_970; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_972 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_1_T_3[5:0] ? buffer_3_9 : _GEN_971; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_973 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_1_T_3[5:0] ? buffer_3_10 : _GEN_972; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_974 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_1_T_3[5:0] ? buffer_3_11 : _GEN_973; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_975 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_1_T_3[5:0] ? buffer_3_12 : _GEN_974; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_976 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_1_T_3[5:0] ? buffer_3_13 : _GEN_975; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_977 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_1_T_3[5:0] ? buffer_3_14 : _GEN_976; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_978 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_1_T_3[5:0] ? buffer_3_15 : _GEN_977; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_979 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_1_T_3[5:0] ? buffer_3_16 : _GEN_978; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_980 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_1_T_3[5:0] ? buffer_3_17 : _GEN_979; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_981 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_1_T_3[5:0] ? buffer_3_18 : _GEN_980; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_982 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_1_T_3[5:0] ? buffer_3_19 : _GEN_981; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_983 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_1_T_3[5:0] ? buffer_3_20 : _GEN_982; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_984 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_1_T_3[5:0] ? buffer_3_21 : _GEN_983; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_985 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_1_T_3[5:0] ? buffer_3_22 : _GEN_984; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_986 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_1_T_3[5:0] ? buffer_3_23 : _GEN_985; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_987 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_1_T_3[5:0] ? buffer_3_24 : _GEN_986; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_988 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_1_T_3[5:0] ? buffer_3_25 : _GEN_987; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_989 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_1_T_3[5:0] ? buffer_3_26 : _GEN_988; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_990 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_1_T_3[5:0] ? buffer_3_27 : _GEN_989; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_991 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_1_T_3[5:0] ? buffer_3_28 : _GEN_990; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_992 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_1_T_3[5:0] ? buffer_3_29 : _GEN_991; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_993 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_1_T_3[5:0] ? buffer_3_30 : _GEN_992; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_994 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_1_T_3[5:0] ? buffer_3_31 : _GEN_993; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_995 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_1_T_3[5:0] ? buffer_3_32 : _GEN_994; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_996 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_1_T_3[5:0] ? buffer_3_33 : _GEN_995; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_997 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_1_T_3[5:0] ? buffer_3_34 : _GEN_996; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_998 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_1_T_3[5:0] ? buffer_3_35 : _GEN_997; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_999 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_1_T_3[5:0] ? buffer_3_36 : _GEN_998; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1000 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_1_T_3[5:0] ? buffer_3_37 : _GEN_999; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1001 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_1_T_3[5:0] ? buffer_3_38 : _GEN_1000; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1002 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_1_T_3[5:0] ? buffer_3_39 : _GEN_1001; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1003 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_1_T_3[5:0] ? buffer_3_40 : _GEN_1002; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1004 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_1_T_3[5:0] ? buffer_3_41 : _GEN_1003; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1005 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_1_T_3[5:0] ? buffer_3_42 : _GEN_1004; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1006 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_1_T_3[5:0] ? buffer_3_43 : _GEN_1005; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1007 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_1_T_3[5:0] ? buffer_3_44 : _GEN_1006; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1008 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_1_T_3[5:0] ? buffer_3_45 : _GEN_1007; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1009 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_1_T_3[5:0] ? buffer_3_46 : _GEN_1008; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1010 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_1_T_3[5:0] ? buffer_3_47 : _GEN_1009; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1011 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_1_T_3[5:0] ? buffer_3_48 : _GEN_1010; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1012 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_1_T_3[5:0] ? buffer_3_49 : _GEN_1011; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1013 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_1_T_3[5:0] ? buffer_3_50 : _GEN_1012; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1014 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_1_T_3[5:0] ? buffer_3_51 : _GEN_1013; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1015 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_1_T_3[5:0] ? buffer_3_52 : _GEN_1014; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1016 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_1_T_3[5:0] ? buffer_3_53 : _GEN_1015; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1017 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_1_T_3[5:0] ? buffer_3_54 : _GEN_1016; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1018 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_1_T_3[5:0] ? buffer_3_55 : _GEN_1017; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1019 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_1_T_3[5:0] ? buffer_3_56 : _GEN_1018; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1020 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_1_T_3[5:0] ? buffer_3_57 : _GEN_1019; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1021 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_1_T_3[5:0] ? buffer_3_58 : _GEN_1020; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1022 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_1_T_3[5:0] ? buffer_3_59 : _GEN_1021; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1023 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_1_T_3[5:0] ? buffer_3_60 : _GEN_1022; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1024 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_1_T_3[5:0] ? buffer_3_61 : _GEN_1023; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1025 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_1_T_3[5:0] ? buffer_3_62 : _GEN_1024; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1026 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_1_T_3[5:0] ? buffer_3_63 : _GEN_1025; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_2_T_3 = _io_out_weight_0_T_1 + 8'h2; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_1028 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_2_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1029 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_2_T_3[5:0] ? buffer_0_2 : _GEN_1028; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1030 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_2_T_3[5:0] ? buffer_0_3 : _GEN_1029; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1031 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_2_T_3[5:0] ? buffer_0_4 : _GEN_1030; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1032 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_2_T_3[5:0] ? buffer_0_5 : _GEN_1031; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1033 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_2_T_3[5:0] ? buffer_0_6 : _GEN_1032; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1034 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_2_T_3[5:0] ? buffer_0_7 : _GEN_1033; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1035 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_2_T_3[5:0] ? buffer_0_8 : _GEN_1034; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1036 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_2_T_3[5:0] ? buffer_0_9 : _GEN_1035; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1037 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_2_T_3[5:0] ? buffer_0_10 : _GEN_1036; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1038 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_2_T_3[5:0] ? buffer_0_11 : _GEN_1037; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1039 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_2_T_3[5:0] ? buffer_0_12 : _GEN_1038; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1040 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_2_T_3[5:0] ? buffer_0_13 : _GEN_1039; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1041 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_2_T_3[5:0] ? buffer_0_14 : _GEN_1040; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1042 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_2_T_3[5:0] ? buffer_0_15 : _GEN_1041; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1043 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_2_T_3[5:0] ? buffer_0_16 : _GEN_1042; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1044 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_2_T_3[5:0] ? buffer_0_17 : _GEN_1043; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1045 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_2_T_3[5:0] ? buffer_0_18 : _GEN_1044; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1046 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_2_T_3[5:0] ? buffer_0_19 : _GEN_1045; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1047 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_2_T_3[5:0] ? buffer_0_20 : _GEN_1046; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1048 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_2_T_3[5:0] ? buffer_0_21 : _GEN_1047; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1049 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_2_T_3[5:0] ? buffer_0_22 : _GEN_1048; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1050 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_2_T_3[5:0] ? buffer_0_23 : _GEN_1049; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1051 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_2_T_3[5:0] ? buffer_0_24 : _GEN_1050; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1052 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_2_T_3[5:0] ? buffer_0_25 : _GEN_1051; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1053 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_2_T_3[5:0] ? buffer_0_26 : _GEN_1052; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1054 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_2_T_3[5:0] ? buffer_0_27 : _GEN_1053; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1055 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_2_T_3[5:0] ? buffer_0_28 : _GEN_1054; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1056 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_2_T_3[5:0] ? buffer_0_29 : _GEN_1055; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1057 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_2_T_3[5:0] ? buffer_0_30 : _GEN_1056; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1058 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_2_T_3[5:0] ? buffer_0_31 : _GEN_1057; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1059 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_2_T_3[5:0] ? buffer_0_32 : _GEN_1058; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1060 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_2_T_3[5:0] ? buffer_0_33 : _GEN_1059; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1061 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_2_T_3[5:0] ? buffer_0_34 : _GEN_1060; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1062 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_2_T_3[5:0] ? buffer_0_35 : _GEN_1061; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1063 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_2_T_3[5:0] ? buffer_0_36 : _GEN_1062; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1064 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_2_T_3[5:0] ? buffer_0_37 : _GEN_1063; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1065 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_2_T_3[5:0] ? buffer_0_38 : _GEN_1064; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1066 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_2_T_3[5:0] ? buffer_0_39 : _GEN_1065; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1067 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_2_T_3[5:0] ? buffer_0_40 : _GEN_1066; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1068 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_2_T_3[5:0] ? buffer_0_41 : _GEN_1067; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1069 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_2_T_3[5:0] ? buffer_0_42 : _GEN_1068; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1070 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_2_T_3[5:0] ? buffer_0_43 : _GEN_1069; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1071 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_2_T_3[5:0] ? buffer_0_44 : _GEN_1070; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1072 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_2_T_3[5:0] ? buffer_0_45 : _GEN_1071; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1073 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_2_T_3[5:0] ? buffer_0_46 : _GEN_1072; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1074 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_2_T_3[5:0] ? buffer_0_47 : _GEN_1073; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1075 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_2_T_3[5:0] ? buffer_0_48 : _GEN_1074; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1076 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_2_T_3[5:0] ? buffer_0_49 : _GEN_1075; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1077 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_2_T_3[5:0] ? buffer_0_50 : _GEN_1076; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1078 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_2_T_3[5:0] ? buffer_0_51 : _GEN_1077; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1079 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_2_T_3[5:0] ? buffer_0_52 : _GEN_1078; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1080 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_2_T_3[5:0] ? buffer_0_53 : _GEN_1079; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1081 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_2_T_3[5:0] ? buffer_0_54 : _GEN_1080; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1082 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_2_T_3[5:0] ? buffer_0_55 : _GEN_1081; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1083 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_2_T_3[5:0] ? buffer_0_56 : _GEN_1082; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1084 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_2_T_3[5:0] ? buffer_0_57 : _GEN_1083; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1085 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_2_T_3[5:0] ? buffer_0_58 : _GEN_1084; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1086 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_2_T_3[5:0] ? buffer_0_59 : _GEN_1085; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1087 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_2_T_3[5:0] ? buffer_0_60 : _GEN_1086; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1088 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_2_T_3[5:0] ? buffer_0_61 : _GEN_1087; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1089 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_2_T_3[5:0] ? buffer_0_62 : _GEN_1088; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1090 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_2_T_3[5:0] ? buffer_0_63 : _GEN_1089; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1091 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_2_T_3[5:0] ? buffer_1_0 : _GEN_1090; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1092 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_2_T_3[5:0] ? buffer_1_1 : _GEN_1091; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1093 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_2_T_3[5:0] ? buffer_1_2 : _GEN_1092; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1094 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_2_T_3[5:0] ? buffer_1_3 : _GEN_1093; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1095 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_2_T_3[5:0] ? buffer_1_4 : _GEN_1094; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1096 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_2_T_3[5:0] ? buffer_1_5 : _GEN_1095; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1097 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_2_T_3[5:0] ? buffer_1_6 : _GEN_1096; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1098 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_2_T_3[5:0] ? buffer_1_7 : _GEN_1097; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1099 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_2_T_3[5:0] ? buffer_1_8 : _GEN_1098; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1100 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_2_T_3[5:0] ? buffer_1_9 : _GEN_1099; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1101 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_2_T_3[5:0] ? buffer_1_10 : _GEN_1100; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1102 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_2_T_3[5:0] ? buffer_1_11 : _GEN_1101; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1103 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_2_T_3[5:0] ? buffer_1_12 : _GEN_1102; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1104 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_2_T_3[5:0] ? buffer_1_13 : _GEN_1103; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1105 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_2_T_3[5:0] ? buffer_1_14 : _GEN_1104; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1106 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_2_T_3[5:0] ? buffer_1_15 : _GEN_1105; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1107 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_2_T_3[5:0] ? buffer_1_16 : _GEN_1106; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1108 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_2_T_3[5:0] ? buffer_1_17 : _GEN_1107; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1109 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_2_T_3[5:0] ? buffer_1_18 : _GEN_1108; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1110 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_2_T_3[5:0] ? buffer_1_19 : _GEN_1109; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1111 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_2_T_3[5:0] ? buffer_1_20 : _GEN_1110; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1112 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_2_T_3[5:0] ? buffer_1_21 : _GEN_1111; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1113 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_2_T_3[5:0] ? buffer_1_22 : _GEN_1112; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1114 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_2_T_3[5:0] ? buffer_1_23 : _GEN_1113; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1115 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_2_T_3[5:0] ? buffer_1_24 : _GEN_1114; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1116 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_2_T_3[5:0] ? buffer_1_25 : _GEN_1115; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1117 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_2_T_3[5:0] ? buffer_1_26 : _GEN_1116; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1118 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_2_T_3[5:0] ? buffer_1_27 : _GEN_1117; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1119 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_2_T_3[5:0] ? buffer_1_28 : _GEN_1118; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1120 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_2_T_3[5:0] ? buffer_1_29 : _GEN_1119; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1121 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_2_T_3[5:0] ? buffer_1_30 : _GEN_1120; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1122 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_2_T_3[5:0] ? buffer_1_31 : _GEN_1121; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1123 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_2_T_3[5:0] ? buffer_1_32 : _GEN_1122; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1124 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_2_T_3[5:0] ? buffer_1_33 : _GEN_1123; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1125 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_2_T_3[5:0] ? buffer_1_34 : _GEN_1124; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1126 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_2_T_3[5:0] ? buffer_1_35 : _GEN_1125; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1127 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_2_T_3[5:0] ? buffer_1_36 : _GEN_1126; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1128 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_2_T_3[5:0] ? buffer_1_37 : _GEN_1127; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1129 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_2_T_3[5:0] ? buffer_1_38 : _GEN_1128; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1130 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_2_T_3[5:0] ? buffer_1_39 : _GEN_1129; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1131 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_2_T_3[5:0] ? buffer_1_40 : _GEN_1130; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1132 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_2_T_3[5:0] ? buffer_1_41 : _GEN_1131; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1133 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_2_T_3[5:0] ? buffer_1_42 : _GEN_1132; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1134 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_2_T_3[5:0] ? buffer_1_43 : _GEN_1133; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1135 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_2_T_3[5:0] ? buffer_1_44 : _GEN_1134; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1136 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_2_T_3[5:0] ? buffer_1_45 : _GEN_1135; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1137 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_2_T_3[5:0] ? buffer_1_46 : _GEN_1136; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1138 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_2_T_3[5:0] ? buffer_1_47 : _GEN_1137; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1139 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_2_T_3[5:0] ? buffer_1_48 : _GEN_1138; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1140 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_2_T_3[5:0] ? buffer_1_49 : _GEN_1139; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1141 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_2_T_3[5:0] ? buffer_1_50 : _GEN_1140; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1142 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_2_T_3[5:0] ? buffer_1_51 : _GEN_1141; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1143 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_2_T_3[5:0] ? buffer_1_52 : _GEN_1142; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1144 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_2_T_3[5:0] ? buffer_1_53 : _GEN_1143; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1145 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_2_T_3[5:0] ? buffer_1_54 : _GEN_1144; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1146 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_2_T_3[5:0] ? buffer_1_55 : _GEN_1145; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1147 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_2_T_3[5:0] ? buffer_1_56 : _GEN_1146; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1148 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_2_T_3[5:0] ? buffer_1_57 : _GEN_1147; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1149 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_2_T_3[5:0] ? buffer_1_58 : _GEN_1148; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1150 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_2_T_3[5:0] ? buffer_1_59 : _GEN_1149; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1151 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_2_T_3[5:0] ? buffer_1_60 : _GEN_1150; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1152 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_2_T_3[5:0] ? buffer_1_61 : _GEN_1151; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1153 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_2_T_3[5:0] ? buffer_1_62 : _GEN_1152; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1154 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_2_T_3[5:0] ? buffer_1_63 : _GEN_1153; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1155 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_2_T_3[5:0] ? buffer_2_0 : _GEN_1154; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1156 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_2_T_3[5:0] ? buffer_2_1 : _GEN_1155; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1157 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_2_T_3[5:0] ? buffer_2_2 : _GEN_1156; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1158 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_2_T_3[5:0] ? buffer_2_3 : _GEN_1157; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1159 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_2_T_3[5:0] ? buffer_2_4 : _GEN_1158; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1160 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_2_T_3[5:0] ? buffer_2_5 : _GEN_1159; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1161 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_2_T_3[5:0] ? buffer_2_6 : _GEN_1160; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1162 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_2_T_3[5:0] ? buffer_2_7 : _GEN_1161; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1163 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_2_T_3[5:0] ? buffer_2_8 : _GEN_1162; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1164 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_2_T_3[5:0] ? buffer_2_9 : _GEN_1163; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1165 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_2_T_3[5:0] ? buffer_2_10 : _GEN_1164; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1166 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_2_T_3[5:0] ? buffer_2_11 : _GEN_1165; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1167 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_2_T_3[5:0] ? buffer_2_12 : _GEN_1166; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1168 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_2_T_3[5:0] ? buffer_2_13 : _GEN_1167; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1169 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_2_T_3[5:0] ? buffer_2_14 : _GEN_1168; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1170 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_2_T_3[5:0] ? buffer_2_15 : _GEN_1169; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1171 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_2_T_3[5:0] ? buffer_2_16 : _GEN_1170; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1172 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_2_T_3[5:0] ? buffer_2_17 : _GEN_1171; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1173 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_2_T_3[5:0] ? buffer_2_18 : _GEN_1172; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1174 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_2_T_3[5:0] ? buffer_2_19 : _GEN_1173; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1175 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_2_T_3[5:0] ? buffer_2_20 : _GEN_1174; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1176 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_2_T_3[5:0] ? buffer_2_21 : _GEN_1175; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1177 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_2_T_3[5:0] ? buffer_2_22 : _GEN_1176; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1178 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_2_T_3[5:0] ? buffer_2_23 : _GEN_1177; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1179 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_2_T_3[5:0] ? buffer_2_24 : _GEN_1178; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1180 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_2_T_3[5:0] ? buffer_2_25 : _GEN_1179; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1181 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_2_T_3[5:0] ? buffer_2_26 : _GEN_1180; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1182 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_2_T_3[5:0] ? buffer_2_27 : _GEN_1181; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1183 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_2_T_3[5:0] ? buffer_2_28 : _GEN_1182; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1184 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_2_T_3[5:0] ? buffer_2_29 : _GEN_1183; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1185 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_2_T_3[5:0] ? buffer_2_30 : _GEN_1184; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1186 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_2_T_3[5:0] ? buffer_2_31 : _GEN_1185; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1187 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_2_T_3[5:0] ? buffer_2_32 : _GEN_1186; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1188 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_2_T_3[5:0] ? buffer_2_33 : _GEN_1187; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1189 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_2_T_3[5:0] ? buffer_2_34 : _GEN_1188; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1190 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_2_T_3[5:0] ? buffer_2_35 : _GEN_1189; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1191 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_2_T_3[5:0] ? buffer_2_36 : _GEN_1190; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1192 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_2_T_3[5:0] ? buffer_2_37 : _GEN_1191; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1193 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_2_T_3[5:0] ? buffer_2_38 : _GEN_1192; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1194 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_2_T_3[5:0] ? buffer_2_39 : _GEN_1193; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1195 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_2_T_3[5:0] ? buffer_2_40 : _GEN_1194; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1196 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_2_T_3[5:0] ? buffer_2_41 : _GEN_1195; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1197 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_2_T_3[5:0] ? buffer_2_42 : _GEN_1196; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1198 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_2_T_3[5:0] ? buffer_2_43 : _GEN_1197; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1199 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_2_T_3[5:0] ? buffer_2_44 : _GEN_1198; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1200 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_2_T_3[5:0] ? buffer_2_45 : _GEN_1199; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1201 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_2_T_3[5:0] ? buffer_2_46 : _GEN_1200; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1202 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_2_T_3[5:0] ? buffer_2_47 : _GEN_1201; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1203 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_2_T_3[5:0] ? buffer_2_48 : _GEN_1202; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1204 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_2_T_3[5:0] ? buffer_2_49 : _GEN_1203; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1205 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_2_T_3[5:0] ? buffer_2_50 : _GEN_1204; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1206 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_2_T_3[5:0] ? buffer_2_51 : _GEN_1205; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1207 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_2_T_3[5:0] ? buffer_2_52 : _GEN_1206; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1208 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_2_T_3[5:0] ? buffer_2_53 : _GEN_1207; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1209 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_2_T_3[5:0] ? buffer_2_54 : _GEN_1208; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1210 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_2_T_3[5:0] ? buffer_2_55 : _GEN_1209; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1211 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_2_T_3[5:0] ? buffer_2_56 : _GEN_1210; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1212 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_2_T_3[5:0] ? buffer_2_57 : _GEN_1211; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1213 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_2_T_3[5:0] ? buffer_2_58 : _GEN_1212; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1214 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_2_T_3[5:0] ? buffer_2_59 : _GEN_1213; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1215 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_2_T_3[5:0] ? buffer_2_60 : _GEN_1214; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1216 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_2_T_3[5:0] ? buffer_2_61 : _GEN_1215; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1217 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_2_T_3[5:0] ? buffer_2_62 : _GEN_1216; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1218 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_2_T_3[5:0] ? buffer_2_63 : _GEN_1217; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1219 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_2_T_3[5:0] ? buffer_3_0 : _GEN_1218; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1220 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_2_T_3[5:0] ? buffer_3_1 : _GEN_1219; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1221 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_2_T_3[5:0] ? buffer_3_2 : _GEN_1220; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1222 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_2_T_3[5:0] ? buffer_3_3 : _GEN_1221; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1223 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_2_T_3[5:0] ? buffer_3_4 : _GEN_1222; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1224 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_2_T_3[5:0] ? buffer_3_5 : _GEN_1223; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1225 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_2_T_3[5:0] ? buffer_3_6 : _GEN_1224; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1226 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_2_T_3[5:0] ? buffer_3_7 : _GEN_1225; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1227 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_2_T_3[5:0] ? buffer_3_8 : _GEN_1226; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1228 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_2_T_3[5:0] ? buffer_3_9 : _GEN_1227; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1229 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_2_T_3[5:0] ? buffer_3_10 : _GEN_1228; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1230 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_2_T_3[5:0] ? buffer_3_11 : _GEN_1229; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1231 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_2_T_3[5:0] ? buffer_3_12 : _GEN_1230; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1232 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_2_T_3[5:0] ? buffer_3_13 : _GEN_1231; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1233 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_2_T_3[5:0] ? buffer_3_14 : _GEN_1232; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1234 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_2_T_3[5:0] ? buffer_3_15 : _GEN_1233; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1235 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_2_T_3[5:0] ? buffer_3_16 : _GEN_1234; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1236 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_2_T_3[5:0] ? buffer_3_17 : _GEN_1235; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1237 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_2_T_3[5:0] ? buffer_3_18 : _GEN_1236; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1238 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_2_T_3[5:0] ? buffer_3_19 : _GEN_1237; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1239 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_2_T_3[5:0] ? buffer_3_20 : _GEN_1238; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1240 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_2_T_3[5:0] ? buffer_3_21 : _GEN_1239; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1241 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_2_T_3[5:0] ? buffer_3_22 : _GEN_1240; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1242 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_2_T_3[5:0] ? buffer_3_23 : _GEN_1241; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1243 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_2_T_3[5:0] ? buffer_3_24 : _GEN_1242; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1244 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_2_T_3[5:0] ? buffer_3_25 : _GEN_1243; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1245 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_2_T_3[5:0] ? buffer_3_26 : _GEN_1244; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1246 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_2_T_3[5:0] ? buffer_3_27 : _GEN_1245; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1247 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_2_T_3[5:0] ? buffer_3_28 : _GEN_1246; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1248 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_2_T_3[5:0] ? buffer_3_29 : _GEN_1247; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1249 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_2_T_3[5:0] ? buffer_3_30 : _GEN_1248; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1250 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_2_T_3[5:0] ? buffer_3_31 : _GEN_1249; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1251 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_2_T_3[5:0] ? buffer_3_32 : _GEN_1250; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1252 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_2_T_3[5:0] ? buffer_3_33 : _GEN_1251; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1253 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_2_T_3[5:0] ? buffer_3_34 : _GEN_1252; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1254 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_2_T_3[5:0] ? buffer_3_35 : _GEN_1253; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1255 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_2_T_3[5:0] ? buffer_3_36 : _GEN_1254; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1256 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_2_T_3[5:0] ? buffer_3_37 : _GEN_1255; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1257 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_2_T_3[5:0] ? buffer_3_38 : _GEN_1256; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1258 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_2_T_3[5:0] ? buffer_3_39 : _GEN_1257; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1259 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_2_T_3[5:0] ? buffer_3_40 : _GEN_1258; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1260 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_2_T_3[5:0] ? buffer_3_41 : _GEN_1259; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1261 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_2_T_3[5:0] ? buffer_3_42 : _GEN_1260; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1262 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_2_T_3[5:0] ? buffer_3_43 : _GEN_1261; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1263 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_2_T_3[5:0] ? buffer_3_44 : _GEN_1262; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1264 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_2_T_3[5:0] ? buffer_3_45 : _GEN_1263; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1265 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_2_T_3[5:0] ? buffer_3_46 : _GEN_1264; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1266 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_2_T_3[5:0] ? buffer_3_47 : _GEN_1265; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1267 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_2_T_3[5:0] ? buffer_3_48 : _GEN_1266; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1268 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_2_T_3[5:0] ? buffer_3_49 : _GEN_1267; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1269 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_2_T_3[5:0] ? buffer_3_50 : _GEN_1268; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1270 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_2_T_3[5:0] ? buffer_3_51 : _GEN_1269; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1271 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_2_T_3[5:0] ? buffer_3_52 : _GEN_1270; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1272 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_2_T_3[5:0] ? buffer_3_53 : _GEN_1271; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1273 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_2_T_3[5:0] ? buffer_3_54 : _GEN_1272; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1274 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_2_T_3[5:0] ? buffer_3_55 : _GEN_1273; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1275 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_2_T_3[5:0] ? buffer_3_56 : _GEN_1274; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1276 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_2_T_3[5:0] ? buffer_3_57 : _GEN_1275; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1277 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_2_T_3[5:0] ? buffer_3_58 : _GEN_1276; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1278 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_2_T_3[5:0] ? buffer_3_59 : _GEN_1277; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1279 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_2_T_3[5:0] ? buffer_3_60 : _GEN_1278; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1280 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_2_T_3[5:0] ? buffer_3_61 : _GEN_1279; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1281 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_2_T_3[5:0] ? buffer_3_62 : _GEN_1280; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1282 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_2_T_3[5:0] ? buffer_3_63 : _GEN_1281; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_3_T_3 = _io_out_weight_0_T_1 + 8'h3; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_1284 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_3_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1285 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_3_T_3[5:0] ? buffer_0_2 : _GEN_1284; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1286 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_3_T_3[5:0] ? buffer_0_3 : _GEN_1285; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1287 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_3_T_3[5:0] ? buffer_0_4 : _GEN_1286; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1288 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_3_T_3[5:0] ? buffer_0_5 : _GEN_1287; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1289 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_3_T_3[5:0] ? buffer_0_6 : _GEN_1288; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1290 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_3_T_3[5:0] ? buffer_0_7 : _GEN_1289; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1291 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_3_T_3[5:0] ? buffer_0_8 : _GEN_1290; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1292 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_3_T_3[5:0] ? buffer_0_9 : _GEN_1291; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1293 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_3_T_3[5:0] ? buffer_0_10 : _GEN_1292; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1294 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_3_T_3[5:0] ? buffer_0_11 : _GEN_1293; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1295 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_3_T_3[5:0] ? buffer_0_12 : _GEN_1294; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1296 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_3_T_3[5:0] ? buffer_0_13 : _GEN_1295; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1297 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_3_T_3[5:0] ? buffer_0_14 : _GEN_1296; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1298 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_3_T_3[5:0] ? buffer_0_15 : _GEN_1297; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1299 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_3_T_3[5:0] ? buffer_0_16 : _GEN_1298; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1300 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_3_T_3[5:0] ? buffer_0_17 : _GEN_1299; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1301 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_3_T_3[5:0] ? buffer_0_18 : _GEN_1300; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1302 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_3_T_3[5:0] ? buffer_0_19 : _GEN_1301; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1303 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_3_T_3[5:0] ? buffer_0_20 : _GEN_1302; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1304 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_3_T_3[5:0] ? buffer_0_21 : _GEN_1303; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1305 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_3_T_3[5:0] ? buffer_0_22 : _GEN_1304; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1306 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_3_T_3[5:0] ? buffer_0_23 : _GEN_1305; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1307 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_3_T_3[5:0] ? buffer_0_24 : _GEN_1306; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1308 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_3_T_3[5:0] ? buffer_0_25 : _GEN_1307; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1309 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_3_T_3[5:0] ? buffer_0_26 : _GEN_1308; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1310 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_3_T_3[5:0] ? buffer_0_27 : _GEN_1309; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1311 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_3_T_3[5:0] ? buffer_0_28 : _GEN_1310; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1312 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_3_T_3[5:0] ? buffer_0_29 : _GEN_1311; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1313 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_3_T_3[5:0] ? buffer_0_30 : _GEN_1312; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1314 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_3_T_3[5:0] ? buffer_0_31 : _GEN_1313; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1315 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_3_T_3[5:0] ? buffer_0_32 : _GEN_1314; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1316 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_3_T_3[5:0] ? buffer_0_33 : _GEN_1315; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1317 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_3_T_3[5:0] ? buffer_0_34 : _GEN_1316; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1318 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_3_T_3[5:0] ? buffer_0_35 : _GEN_1317; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1319 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_3_T_3[5:0] ? buffer_0_36 : _GEN_1318; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1320 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_3_T_3[5:0] ? buffer_0_37 : _GEN_1319; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1321 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_3_T_3[5:0] ? buffer_0_38 : _GEN_1320; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1322 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_3_T_3[5:0] ? buffer_0_39 : _GEN_1321; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1323 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_3_T_3[5:0] ? buffer_0_40 : _GEN_1322; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1324 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_3_T_3[5:0] ? buffer_0_41 : _GEN_1323; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1325 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_3_T_3[5:0] ? buffer_0_42 : _GEN_1324; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1326 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_3_T_3[5:0] ? buffer_0_43 : _GEN_1325; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1327 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_3_T_3[5:0] ? buffer_0_44 : _GEN_1326; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1328 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_3_T_3[5:0] ? buffer_0_45 : _GEN_1327; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1329 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_3_T_3[5:0] ? buffer_0_46 : _GEN_1328; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1330 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_3_T_3[5:0] ? buffer_0_47 : _GEN_1329; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1331 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_3_T_3[5:0] ? buffer_0_48 : _GEN_1330; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1332 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_3_T_3[5:0] ? buffer_0_49 : _GEN_1331; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1333 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_3_T_3[5:0] ? buffer_0_50 : _GEN_1332; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1334 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_3_T_3[5:0] ? buffer_0_51 : _GEN_1333; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1335 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_3_T_3[5:0] ? buffer_0_52 : _GEN_1334; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1336 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_3_T_3[5:0] ? buffer_0_53 : _GEN_1335; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1337 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_3_T_3[5:0] ? buffer_0_54 : _GEN_1336; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1338 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_3_T_3[5:0] ? buffer_0_55 : _GEN_1337; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1339 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_3_T_3[5:0] ? buffer_0_56 : _GEN_1338; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1340 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_3_T_3[5:0] ? buffer_0_57 : _GEN_1339; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1341 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_3_T_3[5:0] ? buffer_0_58 : _GEN_1340; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1342 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_3_T_3[5:0] ? buffer_0_59 : _GEN_1341; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1343 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_3_T_3[5:0] ? buffer_0_60 : _GEN_1342; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1344 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_3_T_3[5:0] ? buffer_0_61 : _GEN_1343; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1345 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_3_T_3[5:0] ? buffer_0_62 : _GEN_1344; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1346 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_3_T_3[5:0] ? buffer_0_63 : _GEN_1345; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1347 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_3_T_3[5:0] ? buffer_1_0 : _GEN_1346; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1348 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_3_T_3[5:0] ? buffer_1_1 : _GEN_1347; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1349 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_3_T_3[5:0] ? buffer_1_2 : _GEN_1348; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1350 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_3_T_3[5:0] ? buffer_1_3 : _GEN_1349; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1351 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_3_T_3[5:0] ? buffer_1_4 : _GEN_1350; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1352 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_3_T_3[5:0] ? buffer_1_5 : _GEN_1351; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1353 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_3_T_3[5:0] ? buffer_1_6 : _GEN_1352; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1354 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_3_T_3[5:0] ? buffer_1_7 : _GEN_1353; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1355 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_3_T_3[5:0] ? buffer_1_8 : _GEN_1354; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1356 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_3_T_3[5:0] ? buffer_1_9 : _GEN_1355; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1357 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_3_T_3[5:0] ? buffer_1_10 : _GEN_1356; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1358 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_3_T_3[5:0] ? buffer_1_11 : _GEN_1357; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1359 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_3_T_3[5:0] ? buffer_1_12 : _GEN_1358; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1360 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_3_T_3[5:0] ? buffer_1_13 : _GEN_1359; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1361 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_3_T_3[5:0] ? buffer_1_14 : _GEN_1360; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1362 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_3_T_3[5:0] ? buffer_1_15 : _GEN_1361; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1363 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_3_T_3[5:0] ? buffer_1_16 : _GEN_1362; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1364 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_3_T_3[5:0] ? buffer_1_17 : _GEN_1363; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1365 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_3_T_3[5:0] ? buffer_1_18 : _GEN_1364; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1366 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_3_T_3[5:0] ? buffer_1_19 : _GEN_1365; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1367 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_3_T_3[5:0] ? buffer_1_20 : _GEN_1366; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1368 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_3_T_3[5:0] ? buffer_1_21 : _GEN_1367; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1369 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_3_T_3[5:0] ? buffer_1_22 : _GEN_1368; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1370 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_3_T_3[5:0] ? buffer_1_23 : _GEN_1369; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1371 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_3_T_3[5:0] ? buffer_1_24 : _GEN_1370; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1372 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_3_T_3[5:0] ? buffer_1_25 : _GEN_1371; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1373 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_3_T_3[5:0] ? buffer_1_26 : _GEN_1372; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1374 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_3_T_3[5:0] ? buffer_1_27 : _GEN_1373; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1375 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_3_T_3[5:0] ? buffer_1_28 : _GEN_1374; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1376 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_3_T_3[5:0] ? buffer_1_29 : _GEN_1375; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1377 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_3_T_3[5:0] ? buffer_1_30 : _GEN_1376; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1378 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_3_T_3[5:0] ? buffer_1_31 : _GEN_1377; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1379 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_3_T_3[5:0] ? buffer_1_32 : _GEN_1378; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1380 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_3_T_3[5:0] ? buffer_1_33 : _GEN_1379; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1381 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_3_T_3[5:0] ? buffer_1_34 : _GEN_1380; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1382 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_3_T_3[5:0] ? buffer_1_35 : _GEN_1381; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1383 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_3_T_3[5:0] ? buffer_1_36 : _GEN_1382; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1384 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_3_T_3[5:0] ? buffer_1_37 : _GEN_1383; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1385 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_3_T_3[5:0] ? buffer_1_38 : _GEN_1384; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1386 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_3_T_3[5:0] ? buffer_1_39 : _GEN_1385; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1387 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_3_T_3[5:0] ? buffer_1_40 : _GEN_1386; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1388 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_3_T_3[5:0] ? buffer_1_41 : _GEN_1387; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1389 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_3_T_3[5:0] ? buffer_1_42 : _GEN_1388; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1390 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_3_T_3[5:0] ? buffer_1_43 : _GEN_1389; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1391 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_3_T_3[5:0] ? buffer_1_44 : _GEN_1390; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1392 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_3_T_3[5:0] ? buffer_1_45 : _GEN_1391; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1393 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_3_T_3[5:0] ? buffer_1_46 : _GEN_1392; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1394 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_3_T_3[5:0] ? buffer_1_47 : _GEN_1393; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1395 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_3_T_3[5:0] ? buffer_1_48 : _GEN_1394; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1396 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_3_T_3[5:0] ? buffer_1_49 : _GEN_1395; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1397 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_3_T_3[5:0] ? buffer_1_50 : _GEN_1396; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1398 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_3_T_3[5:0] ? buffer_1_51 : _GEN_1397; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1399 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_3_T_3[5:0] ? buffer_1_52 : _GEN_1398; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1400 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_3_T_3[5:0] ? buffer_1_53 : _GEN_1399; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1401 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_3_T_3[5:0] ? buffer_1_54 : _GEN_1400; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1402 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_3_T_3[5:0] ? buffer_1_55 : _GEN_1401; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1403 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_3_T_3[5:0] ? buffer_1_56 : _GEN_1402; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1404 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_3_T_3[5:0] ? buffer_1_57 : _GEN_1403; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1405 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_3_T_3[5:0] ? buffer_1_58 : _GEN_1404; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1406 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_3_T_3[5:0] ? buffer_1_59 : _GEN_1405; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1407 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_3_T_3[5:0] ? buffer_1_60 : _GEN_1406; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1408 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_3_T_3[5:0] ? buffer_1_61 : _GEN_1407; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1409 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_3_T_3[5:0] ? buffer_1_62 : _GEN_1408; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1410 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_3_T_3[5:0] ? buffer_1_63 : _GEN_1409; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1411 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_3_T_3[5:0] ? buffer_2_0 : _GEN_1410; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1412 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_3_T_3[5:0] ? buffer_2_1 : _GEN_1411; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1413 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_3_T_3[5:0] ? buffer_2_2 : _GEN_1412; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1414 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_3_T_3[5:0] ? buffer_2_3 : _GEN_1413; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1415 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_3_T_3[5:0] ? buffer_2_4 : _GEN_1414; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1416 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_3_T_3[5:0] ? buffer_2_5 : _GEN_1415; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1417 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_3_T_3[5:0] ? buffer_2_6 : _GEN_1416; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1418 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_3_T_3[5:0] ? buffer_2_7 : _GEN_1417; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1419 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_3_T_3[5:0] ? buffer_2_8 : _GEN_1418; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1420 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_3_T_3[5:0] ? buffer_2_9 : _GEN_1419; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1421 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_3_T_3[5:0] ? buffer_2_10 : _GEN_1420; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1422 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_3_T_3[5:0] ? buffer_2_11 : _GEN_1421; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1423 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_3_T_3[5:0] ? buffer_2_12 : _GEN_1422; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1424 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_3_T_3[5:0] ? buffer_2_13 : _GEN_1423; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1425 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_3_T_3[5:0] ? buffer_2_14 : _GEN_1424; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1426 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_3_T_3[5:0] ? buffer_2_15 : _GEN_1425; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1427 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_3_T_3[5:0] ? buffer_2_16 : _GEN_1426; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1428 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_3_T_3[5:0] ? buffer_2_17 : _GEN_1427; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1429 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_3_T_3[5:0] ? buffer_2_18 : _GEN_1428; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1430 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_3_T_3[5:0] ? buffer_2_19 : _GEN_1429; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1431 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_3_T_3[5:0] ? buffer_2_20 : _GEN_1430; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1432 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_3_T_3[5:0] ? buffer_2_21 : _GEN_1431; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1433 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_3_T_3[5:0] ? buffer_2_22 : _GEN_1432; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1434 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_3_T_3[5:0] ? buffer_2_23 : _GEN_1433; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1435 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_3_T_3[5:0] ? buffer_2_24 : _GEN_1434; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1436 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_3_T_3[5:0] ? buffer_2_25 : _GEN_1435; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1437 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_3_T_3[5:0] ? buffer_2_26 : _GEN_1436; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1438 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_3_T_3[5:0] ? buffer_2_27 : _GEN_1437; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1439 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_3_T_3[5:0] ? buffer_2_28 : _GEN_1438; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1440 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_3_T_3[5:0] ? buffer_2_29 : _GEN_1439; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1441 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_3_T_3[5:0] ? buffer_2_30 : _GEN_1440; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1442 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_3_T_3[5:0] ? buffer_2_31 : _GEN_1441; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1443 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_3_T_3[5:0] ? buffer_2_32 : _GEN_1442; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1444 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_3_T_3[5:0] ? buffer_2_33 : _GEN_1443; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1445 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_3_T_3[5:0] ? buffer_2_34 : _GEN_1444; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1446 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_3_T_3[5:0] ? buffer_2_35 : _GEN_1445; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1447 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_3_T_3[5:0] ? buffer_2_36 : _GEN_1446; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1448 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_3_T_3[5:0] ? buffer_2_37 : _GEN_1447; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1449 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_3_T_3[5:0] ? buffer_2_38 : _GEN_1448; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1450 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_3_T_3[5:0] ? buffer_2_39 : _GEN_1449; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1451 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_3_T_3[5:0] ? buffer_2_40 : _GEN_1450; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1452 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_3_T_3[5:0] ? buffer_2_41 : _GEN_1451; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1453 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_3_T_3[5:0] ? buffer_2_42 : _GEN_1452; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1454 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_3_T_3[5:0] ? buffer_2_43 : _GEN_1453; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1455 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_3_T_3[5:0] ? buffer_2_44 : _GEN_1454; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1456 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_3_T_3[5:0] ? buffer_2_45 : _GEN_1455; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1457 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_3_T_3[5:0] ? buffer_2_46 : _GEN_1456; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1458 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_3_T_3[5:0] ? buffer_2_47 : _GEN_1457; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1459 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_3_T_3[5:0] ? buffer_2_48 : _GEN_1458; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1460 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_3_T_3[5:0] ? buffer_2_49 : _GEN_1459; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1461 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_3_T_3[5:0] ? buffer_2_50 : _GEN_1460; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1462 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_3_T_3[5:0] ? buffer_2_51 : _GEN_1461; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1463 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_3_T_3[5:0] ? buffer_2_52 : _GEN_1462; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1464 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_3_T_3[5:0] ? buffer_2_53 : _GEN_1463; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1465 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_3_T_3[5:0] ? buffer_2_54 : _GEN_1464; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1466 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_3_T_3[5:0] ? buffer_2_55 : _GEN_1465; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1467 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_3_T_3[5:0] ? buffer_2_56 : _GEN_1466; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1468 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_3_T_3[5:0] ? buffer_2_57 : _GEN_1467; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1469 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_3_T_3[5:0] ? buffer_2_58 : _GEN_1468; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1470 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_3_T_3[5:0] ? buffer_2_59 : _GEN_1469; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1471 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_3_T_3[5:0] ? buffer_2_60 : _GEN_1470; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1472 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_3_T_3[5:0] ? buffer_2_61 : _GEN_1471; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1473 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_3_T_3[5:0] ? buffer_2_62 : _GEN_1472; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1474 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_3_T_3[5:0] ? buffer_2_63 : _GEN_1473; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1475 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_3_T_3[5:0] ? buffer_3_0 : _GEN_1474; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1476 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_3_T_3[5:0] ? buffer_3_1 : _GEN_1475; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1477 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_3_T_3[5:0] ? buffer_3_2 : _GEN_1476; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1478 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_3_T_3[5:0] ? buffer_3_3 : _GEN_1477; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1479 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_3_T_3[5:0] ? buffer_3_4 : _GEN_1478; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1480 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_3_T_3[5:0] ? buffer_3_5 : _GEN_1479; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1481 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_3_T_3[5:0] ? buffer_3_6 : _GEN_1480; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1482 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_3_T_3[5:0] ? buffer_3_7 : _GEN_1481; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1483 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_3_T_3[5:0] ? buffer_3_8 : _GEN_1482; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1484 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_3_T_3[5:0] ? buffer_3_9 : _GEN_1483; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1485 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_3_T_3[5:0] ? buffer_3_10 : _GEN_1484; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1486 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_3_T_3[5:0] ? buffer_3_11 : _GEN_1485; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1487 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_3_T_3[5:0] ? buffer_3_12 : _GEN_1486; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1488 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_3_T_3[5:0] ? buffer_3_13 : _GEN_1487; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1489 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_3_T_3[5:0] ? buffer_3_14 : _GEN_1488; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1490 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_3_T_3[5:0] ? buffer_3_15 : _GEN_1489; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1491 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_3_T_3[5:0] ? buffer_3_16 : _GEN_1490; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1492 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_3_T_3[5:0] ? buffer_3_17 : _GEN_1491; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1493 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_3_T_3[5:0] ? buffer_3_18 : _GEN_1492; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1494 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_3_T_3[5:0] ? buffer_3_19 : _GEN_1493; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1495 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_3_T_3[5:0] ? buffer_3_20 : _GEN_1494; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1496 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_3_T_3[5:0] ? buffer_3_21 : _GEN_1495; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1497 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_3_T_3[5:0] ? buffer_3_22 : _GEN_1496; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1498 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_3_T_3[5:0] ? buffer_3_23 : _GEN_1497; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1499 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_3_T_3[5:0] ? buffer_3_24 : _GEN_1498; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1500 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_3_T_3[5:0] ? buffer_3_25 : _GEN_1499; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1501 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_3_T_3[5:0] ? buffer_3_26 : _GEN_1500; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1502 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_3_T_3[5:0] ? buffer_3_27 : _GEN_1501; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1503 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_3_T_3[5:0] ? buffer_3_28 : _GEN_1502; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1504 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_3_T_3[5:0] ? buffer_3_29 : _GEN_1503; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1505 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_3_T_3[5:0] ? buffer_3_30 : _GEN_1504; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1506 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_3_T_3[5:0] ? buffer_3_31 : _GEN_1505; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1507 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_3_T_3[5:0] ? buffer_3_32 : _GEN_1506; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1508 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_3_T_3[5:0] ? buffer_3_33 : _GEN_1507; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1509 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_3_T_3[5:0] ? buffer_3_34 : _GEN_1508; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1510 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_3_T_3[5:0] ? buffer_3_35 : _GEN_1509; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1511 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_3_T_3[5:0] ? buffer_3_36 : _GEN_1510; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1512 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_3_T_3[5:0] ? buffer_3_37 : _GEN_1511; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1513 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_3_T_3[5:0] ? buffer_3_38 : _GEN_1512; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1514 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_3_T_3[5:0] ? buffer_3_39 : _GEN_1513; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1515 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_3_T_3[5:0] ? buffer_3_40 : _GEN_1514; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1516 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_3_T_3[5:0] ? buffer_3_41 : _GEN_1515; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1517 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_3_T_3[5:0] ? buffer_3_42 : _GEN_1516; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1518 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_3_T_3[5:0] ? buffer_3_43 : _GEN_1517; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1519 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_3_T_3[5:0] ? buffer_3_44 : _GEN_1518; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1520 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_3_T_3[5:0] ? buffer_3_45 : _GEN_1519; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1521 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_3_T_3[5:0] ? buffer_3_46 : _GEN_1520; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1522 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_3_T_3[5:0] ? buffer_3_47 : _GEN_1521; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1523 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_3_T_3[5:0] ? buffer_3_48 : _GEN_1522; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1524 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_3_T_3[5:0] ? buffer_3_49 : _GEN_1523; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1525 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_3_T_3[5:0] ? buffer_3_50 : _GEN_1524; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1526 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_3_T_3[5:0] ? buffer_3_51 : _GEN_1525; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1527 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_3_T_3[5:0] ? buffer_3_52 : _GEN_1526; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1528 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_3_T_3[5:0] ? buffer_3_53 : _GEN_1527; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1529 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_3_T_3[5:0] ? buffer_3_54 : _GEN_1528; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1530 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_3_T_3[5:0] ? buffer_3_55 : _GEN_1529; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1531 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_3_T_3[5:0] ? buffer_3_56 : _GEN_1530; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1532 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_3_T_3[5:0] ? buffer_3_57 : _GEN_1531; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1533 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_3_T_3[5:0] ? buffer_3_58 : _GEN_1532; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1534 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_3_T_3[5:0] ? buffer_3_59 : _GEN_1533; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1535 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_3_T_3[5:0] ? buffer_3_60 : _GEN_1534; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1536 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_3_T_3[5:0] ? buffer_3_61 : _GEN_1535; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1537 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_3_T_3[5:0] ? buffer_3_62 : _GEN_1536; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1538 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_3_T_3[5:0] ? buffer_3_63 : _GEN_1537; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_4_T_3 = _io_out_weight_0_T_1 + 8'h4; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_1540 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_4_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1541 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_4_T_3[5:0] ? buffer_0_2 : _GEN_1540; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1542 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_4_T_3[5:0] ? buffer_0_3 : _GEN_1541; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1543 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_4_T_3[5:0] ? buffer_0_4 : _GEN_1542; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1544 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_4_T_3[5:0] ? buffer_0_5 : _GEN_1543; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1545 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_4_T_3[5:0] ? buffer_0_6 : _GEN_1544; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1546 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_4_T_3[5:0] ? buffer_0_7 : _GEN_1545; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1547 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_4_T_3[5:0] ? buffer_0_8 : _GEN_1546; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1548 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_4_T_3[5:0] ? buffer_0_9 : _GEN_1547; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1549 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_4_T_3[5:0] ? buffer_0_10 : _GEN_1548; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1550 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_4_T_3[5:0] ? buffer_0_11 : _GEN_1549; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1551 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_4_T_3[5:0] ? buffer_0_12 : _GEN_1550; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1552 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_4_T_3[5:0] ? buffer_0_13 : _GEN_1551; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1553 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_4_T_3[5:0] ? buffer_0_14 : _GEN_1552; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1554 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_4_T_3[5:0] ? buffer_0_15 : _GEN_1553; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1555 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_4_T_3[5:0] ? buffer_0_16 : _GEN_1554; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1556 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_4_T_3[5:0] ? buffer_0_17 : _GEN_1555; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1557 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_4_T_3[5:0] ? buffer_0_18 : _GEN_1556; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1558 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_4_T_3[5:0] ? buffer_0_19 : _GEN_1557; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1559 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_4_T_3[5:0] ? buffer_0_20 : _GEN_1558; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1560 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_4_T_3[5:0] ? buffer_0_21 : _GEN_1559; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1561 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_4_T_3[5:0] ? buffer_0_22 : _GEN_1560; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1562 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_4_T_3[5:0] ? buffer_0_23 : _GEN_1561; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1563 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_4_T_3[5:0] ? buffer_0_24 : _GEN_1562; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1564 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_4_T_3[5:0] ? buffer_0_25 : _GEN_1563; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1565 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_4_T_3[5:0] ? buffer_0_26 : _GEN_1564; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1566 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_4_T_3[5:0] ? buffer_0_27 : _GEN_1565; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1567 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_4_T_3[5:0] ? buffer_0_28 : _GEN_1566; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1568 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_4_T_3[5:0] ? buffer_0_29 : _GEN_1567; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1569 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_4_T_3[5:0] ? buffer_0_30 : _GEN_1568; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1570 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_4_T_3[5:0] ? buffer_0_31 : _GEN_1569; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1571 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_4_T_3[5:0] ? buffer_0_32 : _GEN_1570; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1572 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_4_T_3[5:0] ? buffer_0_33 : _GEN_1571; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1573 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_4_T_3[5:0] ? buffer_0_34 : _GEN_1572; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1574 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_4_T_3[5:0] ? buffer_0_35 : _GEN_1573; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1575 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_4_T_3[5:0] ? buffer_0_36 : _GEN_1574; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1576 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_4_T_3[5:0] ? buffer_0_37 : _GEN_1575; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1577 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_4_T_3[5:0] ? buffer_0_38 : _GEN_1576; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1578 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_4_T_3[5:0] ? buffer_0_39 : _GEN_1577; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1579 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_4_T_3[5:0] ? buffer_0_40 : _GEN_1578; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1580 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_4_T_3[5:0] ? buffer_0_41 : _GEN_1579; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1581 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_4_T_3[5:0] ? buffer_0_42 : _GEN_1580; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1582 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_4_T_3[5:0] ? buffer_0_43 : _GEN_1581; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1583 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_4_T_3[5:0] ? buffer_0_44 : _GEN_1582; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1584 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_4_T_3[5:0] ? buffer_0_45 : _GEN_1583; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1585 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_4_T_3[5:0] ? buffer_0_46 : _GEN_1584; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1586 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_4_T_3[5:0] ? buffer_0_47 : _GEN_1585; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1587 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_4_T_3[5:0] ? buffer_0_48 : _GEN_1586; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1588 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_4_T_3[5:0] ? buffer_0_49 : _GEN_1587; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1589 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_4_T_3[5:0] ? buffer_0_50 : _GEN_1588; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1590 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_4_T_3[5:0] ? buffer_0_51 : _GEN_1589; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1591 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_4_T_3[5:0] ? buffer_0_52 : _GEN_1590; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1592 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_4_T_3[5:0] ? buffer_0_53 : _GEN_1591; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1593 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_4_T_3[5:0] ? buffer_0_54 : _GEN_1592; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1594 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_4_T_3[5:0] ? buffer_0_55 : _GEN_1593; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1595 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_4_T_3[5:0] ? buffer_0_56 : _GEN_1594; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1596 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_4_T_3[5:0] ? buffer_0_57 : _GEN_1595; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1597 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_4_T_3[5:0] ? buffer_0_58 : _GEN_1596; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1598 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_4_T_3[5:0] ? buffer_0_59 : _GEN_1597; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1599 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_4_T_3[5:0] ? buffer_0_60 : _GEN_1598; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1600 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_4_T_3[5:0] ? buffer_0_61 : _GEN_1599; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1601 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_4_T_3[5:0] ? buffer_0_62 : _GEN_1600; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1602 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_4_T_3[5:0] ? buffer_0_63 : _GEN_1601; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1603 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_4_T_3[5:0] ? buffer_1_0 : _GEN_1602; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1604 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_4_T_3[5:0] ? buffer_1_1 : _GEN_1603; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1605 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_4_T_3[5:0] ? buffer_1_2 : _GEN_1604; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1606 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_4_T_3[5:0] ? buffer_1_3 : _GEN_1605; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1607 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_4_T_3[5:0] ? buffer_1_4 : _GEN_1606; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1608 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_4_T_3[5:0] ? buffer_1_5 : _GEN_1607; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1609 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_4_T_3[5:0] ? buffer_1_6 : _GEN_1608; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1610 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_4_T_3[5:0] ? buffer_1_7 : _GEN_1609; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1611 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_4_T_3[5:0] ? buffer_1_8 : _GEN_1610; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1612 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_4_T_3[5:0] ? buffer_1_9 : _GEN_1611; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1613 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_4_T_3[5:0] ? buffer_1_10 : _GEN_1612; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1614 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_4_T_3[5:0] ? buffer_1_11 : _GEN_1613; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1615 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_4_T_3[5:0] ? buffer_1_12 : _GEN_1614; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1616 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_4_T_3[5:0] ? buffer_1_13 : _GEN_1615; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1617 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_4_T_3[5:0] ? buffer_1_14 : _GEN_1616; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1618 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_4_T_3[5:0] ? buffer_1_15 : _GEN_1617; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1619 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_4_T_3[5:0] ? buffer_1_16 : _GEN_1618; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1620 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_4_T_3[5:0] ? buffer_1_17 : _GEN_1619; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1621 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_4_T_3[5:0] ? buffer_1_18 : _GEN_1620; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1622 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_4_T_3[5:0] ? buffer_1_19 : _GEN_1621; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1623 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_4_T_3[5:0] ? buffer_1_20 : _GEN_1622; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1624 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_4_T_3[5:0] ? buffer_1_21 : _GEN_1623; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1625 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_4_T_3[5:0] ? buffer_1_22 : _GEN_1624; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1626 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_4_T_3[5:0] ? buffer_1_23 : _GEN_1625; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1627 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_4_T_3[5:0] ? buffer_1_24 : _GEN_1626; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1628 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_4_T_3[5:0] ? buffer_1_25 : _GEN_1627; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1629 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_4_T_3[5:0] ? buffer_1_26 : _GEN_1628; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1630 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_4_T_3[5:0] ? buffer_1_27 : _GEN_1629; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1631 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_4_T_3[5:0] ? buffer_1_28 : _GEN_1630; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1632 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_4_T_3[5:0] ? buffer_1_29 : _GEN_1631; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1633 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_4_T_3[5:0] ? buffer_1_30 : _GEN_1632; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1634 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_4_T_3[5:0] ? buffer_1_31 : _GEN_1633; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1635 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_4_T_3[5:0] ? buffer_1_32 : _GEN_1634; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1636 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_4_T_3[5:0] ? buffer_1_33 : _GEN_1635; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1637 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_4_T_3[5:0] ? buffer_1_34 : _GEN_1636; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1638 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_4_T_3[5:0] ? buffer_1_35 : _GEN_1637; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1639 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_4_T_3[5:0] ? buffer_1_36 : _GEN_1638; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1640 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_4_T_3[5:0] ? buffer_1_37 : _GEN_1639; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1641 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_4_T_3[5:0] ? buffer_1_38 : _GEN_1640; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1642 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_4_T_3[5:0] ? buffer_1_39 : _GEN_1641; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1643 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_4_T_3[5:0] ? buffer_1_40 : _GEN_1642; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1644 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_4_T_3[5:0] ? buffer_1_41 : _GEN_1643; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1645 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_4_T_3[5:0] ? buffer_1_42 : _GEN_1644; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1646 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_4_T_3[5:0] ? buffer_1_43 : _GEN_1645; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1647 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_4_T_3[5:0] ? buffer_1_44 : _GEN_1646; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1648 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_4_T_3[5:0] ? buffer_1_45 : _GEN_1647; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1649 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_4_T_3[5:0] ? buffer_1_46 : _GEN_1648; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1650 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_4_T_3[5:0] ? buffer_1_47 : _GEN_1649; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1651 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_4_T_3[5:0] ? buffer_1_48 : _GEN_1650; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1652 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_4_T_3[5:0] ? buffer_1_49 : _GEN_1651; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1653 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_4_T_3[5:0] ? buffer_1_50 : _GEN_1652; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1654 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_4_T_3[5:0] ? buffer_1_51 : _GEN_1653; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1655 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_4_T_3[5:0] ? buffer_1_52 : _GEN_1654; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1656 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_4_T_3[5:0] ? buffer_1_53 : _GEN_1655; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1657 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_4_T_3[5:0] ? buffer_1_54 : _GEN_1656; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1658 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_4_T_3[5:0] ? buffer_1_55 : _GEN_1657; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1659 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_4_T_3[5:0] ? buffer_1_56 : _GEN_1658; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1660 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_4_T_3[5:0] ? buffer_1_57 : _GEN_1659; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1661 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_4_T_3[5:0] ? buffer_1_58 : _GEN_1660; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1662 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_4_T_3[5:0] ? buffer_1_59 : _GEN_1661; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1663 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_4_T_3[5:0] ? buffer_1_60 : _GEN_1662; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1664 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_4_T_3[5:0] ? buffer_1_61 : _GEN_1663; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1665 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_4_T_3[5:0] ? buffer_1_62 : _GEN_1664; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1666 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_4_T_3[5:0] ? buffer_1_63 : _GEN_1665; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1667 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_4_T_3[5:0] ? buffer_2_0 : _GEN_1666; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1668 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_4_T_3[5:0] ? buffer_2_1 : _GEN_1667; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1669 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_4_T_3[5:0] ? buffer_2_2 : _GEN_1668; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1670 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_4_T_3[5:0] ? buffer_2_3 : _GEN_1669; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1671 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_4_T_3[5:0] ? buffer_2_4 : _GEN_1670; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1672 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_4_T_3[5:0] ? buffer_2_5 : _GEN_1671; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1673 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_4_T_3[5:0] ? buffer_2_6 : _GEN_1672; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1674 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_4_T_3[5:0] ? buffer_2_7 : _GEN_1673; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1675 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_4_T_3[5:0] ? buffer_2_8 : _GEN_1674; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1676 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_4_T_3[5:0] ? buffer_2_9 : _GEN_1675; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1677 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_4_T_3[5:0] ? buffer_2_10 : _GEN_1676; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1678 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_4_T_3[5:0] ? buffer_2_11 : _GEN_1677; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1679 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_4_T_3[5:0] ? buffer_2_12 : _GEN_1678; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1680 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_4_T_3[5:0] ? buffer_2_13 : _GEN_1679; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1681 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_4_T_3[5:0] ? buffer_2_14 : _GEN_1680; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1682 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_4_T_3[5:0] ? buffer_2_15 : _GEN_1681; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1683 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_4_T_3[5:0] ? buffer_2_16 : _GEN_1682; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1684 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_4_T_3[5:0] ? buffer_2_17 : _GEN_1683; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1685 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_4_T_3[5:0] ? buffer_2_18 : _GEN_1684; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1686 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_4_T_3[5:0] ? buffer_2_19 : _GEN_1685; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1687 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_4_T_3[5:0] ? buffer_2_20 : _GEN_1686; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1688 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_4_T_3[5:0] ? buffer_2_21 : _GEN_1687; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1689 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_4_T_3[5:0] ? buffer_2_22 : _GEN_1688; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1690 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_4_T_3[5:0] ? buffer_2_23 : _GEN_1689; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1691 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_4_T_3[5:0] ? buffer_2_24 : _GEN_1690; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1692 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_4_T_3[5:0] ? buffer_2_25 : _GEN_1691; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1693 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_4_T_3[5:0] ? buffer_2_26 : _GEN_1692; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1694 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_4_T_3[5:0] ? buffer_2_27 : _GEN_1693; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1695 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_4_T_3[5:0] ? buffer_2_28 : _GEN_1694; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1696 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_4_T_3[5:0] ? buffer_2_29 : _GEN_1695; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1697 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_4_T_3[5:0] ? buffer_2_30 : _GEN_1696; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1698 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_4_T_3[5:0] ? buffer_2_31 : _GEN_1697; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1699 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_4_T_3[5:0] ? buffer_2_32 : _GEN_1698; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1700 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_4_T_3[5:0] ? buffer_2_33 : _GEN_1699; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1701 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_4_T_3[5:0] ? buffer_2_34 : _GEN_1700; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1702 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_4_T_3[5:0] ? buffer_2_35 : _GEN_1701; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1703 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_4_T_3[5:0] ? buffer_2_36 : _GEN_1702; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1704 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_4_T_3[5:0] ? buffer_2_37 : _GEN_1703; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1705 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_4_T_3[5:0] ? buffer_2_38 : _GEN_1704; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1706 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_4_T_3[5:0] ? buffer_2_39 : _GEN_1705; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1707 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_4_T_3[5:0] ? buffer_2_40 : _GEN_1706; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1708 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_4_T_3[5:0] ? buffer_2_41 : _GEN_1707; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1709 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_4_T_3[5:0] ? buffer_2_42 : _GEN_1708; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1710 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_4_T_3[5:0] ? buffer_2_43 : _GEN_1709; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1711 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_4_T_3[5:0] ? buffer_2_44 : _GEN_1710; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1712 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_4_T_3[5:0] ? buffer_2_45 : _GEN_1711; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1713 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_4_T_3[5:0] ? buffer_2_46 : _GEN_1712; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1714 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_4_T_3[5:0] ? buffer_2_47 : _GEN_1713; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1715 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_4_T_3[5:0] ? buffer_2_48 : _GEN_1714; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1716 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_4_T_3[5:0] ? buffer_2_49 : _GEN_1715; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1717 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_4_T_3[5:0] ? buffer_2_50 : _GEN_1716; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1718 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_4_T_3[5:0] ? buffer_2_51 : _GEN_1717; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1719 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_4_T_3[5:0] ? buffer_2_52 : _GEN_1718; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1720 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_4_T_3[5:0] ? buffer_2_53 : _GEN_1719; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1721 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_4_T_3[5:0] ? buffer_2_54 : _GEN_1720; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1722 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_4_T_3[5:0] ? buffer_2_55 : _GEN_1721; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1723 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_4_T_3[5:0] ? buffer_2_56 : _GEN_1722; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1724 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_4_T_3[5:0] ? buffer_2_57 : _GEN_1723; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1725 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_4_T_3[5:0] ? buffer_2_58 : _GEN_1724; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1726 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_4_T_3[5:0] ? buffer_2_59 : _GEN_1725; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1727 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_4_T_3[5:0] ? buffer_2_60 : _GEN_1726; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1728 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_4_T_3[5:0] ? buffer_2_61 : _GEN_1727; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1729 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_4_T_3[5:0] ? buffer_2_62 : _GEN_1728; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1730 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_4_T_3[5:0] ? buffer_2_63 : _GEN_1729; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1731 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_4_T_3[5:0] ? buffer_3_0 : _GEN_1730; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1732 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_4_T_3[5:0] ? buffer_3_1 : _GEN_1731; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1733 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_4_T_3[5:0] ? buffer_3_2 : _GEN_1732; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1734 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_4_T_3[5:0] ? buffer_3_3 : _GEN_1733; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1735 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_4_T_3[5:0] ? buffer_3_4 : _GEN_1734; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1736 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_4_T_3[5:0] ? buffer_3_5 : _GEN_1735; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1737 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_4_T_3[5:0] ? buffer_3_6 : _GEN_1736; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1738 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_4_T_3[5:0] ? buffer_3_7 : _GEN_1737; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1739 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_4_T_3[5:0] ? buffer_3_8 : _GEN_1738; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1740 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_4_T_3[5:0] ? buffer_3_9 : _GEN_1739; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1741 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_4_T_3[5:0] ? buffer_3_10 : _GEN_1740; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1742 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_4_T_3[5:0] ? buffer_3_11 : _GEN_1741; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1743 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_4_T_3[5:0] ? buffer_3_12 : _GEN_1742; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1744 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_4_T_3[5:0] ? buffer_3_13 : _GEN_1743; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1745 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_4_T_3[5:0] ? buffer_3_14 : _GEN_1744; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1746 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_4_T_3[5:0] ? buffer_3_15 : _GEN_1745; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1747 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_4_T_3[5:0] ? buffer_3_16 : _GEN_1746; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1748 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_4_T_3[5:0] ? buffer_3_17 : _GEN_1747; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1749 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_4_T_3[5:0] ? buffer_3_18 : _GEN_1748; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1750 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_4_T_3[5:0] ? buffer_3_19 : _GEN_1749; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1751 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_4_T_3[5:0] ? buffer_3_20 : _GEN_1750; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1752 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_4_T_3[5:0] ? buffer_3_21 : _GEN_1751; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1753 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_4_T_3[5:0] ? buffer_3_22 : _GEN_1752; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1754 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_4_T_3[5:0] ? buffer_3_23 : _GEN_1753; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1755 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_4_T_3[5:0] ? buffer_3_24 : _GEN_1754; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1756 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_4_T_3[5:0] ? buffer_3_25 : _GEN_1755; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1757 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_4_T_3[5:0] ? buffer_3_26 : _GEN_1756; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1758 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_4_T_3[5:0] ? buffer_3_27 : _GEN_1757; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1759 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_4_T_3[5:0] ? buffer_3_28 : _GEN_1758; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1760 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_4_T_3[5:0] ? buffer_3_29 : _GEN_1759; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1761 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_4_T_3[5:0] ? buffer_3_30 : _GEN_1760; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1762 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_4_T_3[5:0] ? buffer_3_31 : _GEN_1761; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1763 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_4_T_3[5:0] ? buffer_3_32 : _GEN_1762; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1764 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_4_T_3[5:0] ? buffer_3_33 : _GEN_1763; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1765 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_4_T_3[5:0] ? buffer_3_34 : _GEN_1764; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1766 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_4_T_3[5:0] ? buffer_3_35 : _GEN_1765; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1767 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_4_T_3[5:0] ? buffer_3_36 : _GEN_1766; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1768 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_4_T_3[5:0] ? buffer_3_37 : _GEN_1767; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1769 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_4_T_3[5:0] ? buffer_3_38 : _GEN_1768; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1770 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_4_T_3[5:0] ? buffer_3_39 : _GEN_1769; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1771 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_4_T_3[5:0] ? buffer_3_40 : _GEN_1770; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1772 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_4_T_3[5:0] ? buffer_3_41 : _GEN_1771; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1773 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_4_T_3[5:0] ? buffer_3_42 : _GEN_1772; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1774 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_4_T_3[5:0] ? buffer_3_43 : _GEN_1773; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1775 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_4_T_3[5:0] ? buffer_3_44 : _GEN_1774; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1776 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_4_T_3[5:0] ? buffer_3_45 : _GEN_1775; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1777 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_4_T_3[5:0] ? buffer_3_46 : _GEN_1776; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1778 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_4_T_3[5:0] ? buffer_3_47 : _GEN_1777; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1779 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_4_T_3[5:0] ? buffer_3_48 : _GEN_1778; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1780 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_4_T_3[5:0] ? buffer_3_49 : _GEN_1779; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1781 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_4_T_3[5:0] ? buffer_3_50 : _GEN_1780; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1782 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_4_T_3[5:0] ? buffer_3_51 : _GEN_1781; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1783 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_4_T_3[5:0] ? buffer_3_52 : _GEN_1782; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1784 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_4_T_3[5:0] ? buffer_3_53 : _GEN_1783; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1785 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_4_T_3[5:0] ? buffer_3_54 : _GEN_1784; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1786 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_4_T_3[5:0] ? buffer_3_55 : _GEN_1785; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1787 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_4_T_3[5:0] ? buffer_3_56 : _GEN_1786; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1788 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_4_T_3[5:0] ? buffer_3_57 : _GEN_1787; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1789 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_4_T_3[5:0] ? buffer_3_58 : _GEN_1788; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1790 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_4_T_3[5:0] ? buffer_3_59 : _GEN_1789; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1791 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_4_T_3[5:0] ? buffer_3_60 : _GEN_1790; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1792 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_4_T_3[5:0] ? buffer_3_61 : _GEN_1791; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1793 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_4_T_3[5:0] ? buffer_3_62 : _GEN_1792; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1794 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_4_T_3[5:0] ? buffer_3_63 : _GEN_1793; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_5_T_3 = _io_out_weight_0_T_1 + 8'h5; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_1796 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_5_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1797 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_5_T_3[5:0] ? buffer_0_2 : _GEN_1796; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1798 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_5_T_3[5:0] ? buffer_0_3 : _GEN_1797; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1799 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_5_T_3[5:0] ? buffer_0_4 : _GEN_1798; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1800 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_5_T_3[5:0] ? buffer_0_5 : _GEN_1799; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1801 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_5_T_3[5:0] ? buffer_0_6 : _GEN_1800; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1802 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_5_T_3[5:0] ? buffer_0_7 : _GEN_1801; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1803 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_5_T_3[5:0] ? buffer_0_8 : _GEN_1802; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1804 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_5_T_3[5:0] ? buffer_0_9 : _GEN_1803; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1805 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_5_T_3[5:0] ? buffer_0_10 : _GEN_1804; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1806 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_5_T_3[5:0] ? buffer_0_11 : _GEN_1805; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1807 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_5_T_3[5:0] ? buffer_0_12 : _GEN_1806; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1808 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_5_T_3[5:0] ? buffer_0_13 : _GEN_1807; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1809 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_5_T_3[5:0] ? buffer_0_14 : _GEN_1808; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1810 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_5_T_3[5:0] ? buffer_0_15 : _GEN_1809; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1811 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_5_T_3[5:0] ? buffer_0_16 : _GEN_1810; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1812 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_5_T_3[5:0] ? buffer_0_17 : _GEN_1811; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1813 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_5_T_3[5:0] ? buffer_0_18 : _GEN_1812; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1814 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_5_T_3[5:0] ? buffer_0_19 : _GEN_1813; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1815 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_5_T_3[5:0] ? buffer_0_20 : _GEN_1814; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1816 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_5_T_3[5:0] ? buffer_0_21 : _GEN_1815; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1817 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_5_T_3[5:0] ? buffer_0_22 : _GEN_1816; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1818 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_5_T_3[5:0] ? buffer_0_23 : _GEN_1817; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1819 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_5_T_3[5:0] ? buffer_0_24 : _GEN_1818; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1820 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_5_T_3[5:0] ? buffer_0_25 : _GEN_1819; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1821 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_5_T_3[5:0] ? buffer_0_26 : _GEN_1820; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1822 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_5_T_3[5:0] ? buffer_0_27 : _GEN_1821; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1823 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_5_T_3[5:0] ? buffer_0_28 : _GEN_1822; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1824 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_5_T_3[5:0] ? buffer_0_29 : _GEN_1823; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1825 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_5_T_3[5:0] ? buffer_0_30 : _GEN_1824; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1826 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_5_T_3[5:0] ? buffer_0_31 : _GEN_1825; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1827 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_5_T_3[5:0] ? buffer_0_32 : _GEN_1826; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1828 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_5_T_3[5:0] ? buffer_0_33 : _GEN_1827; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1829 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_5_T_3[5:0] ? buffer_0_34 : _GEN_1828; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1830 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_5_T_3[5:0] ? buffer_0_35 : _GEN_1829; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1831 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_5_T_3[5:0] ? buffer_0_36 : _GEN_1830; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1832 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_5_T_3[5:0] ? buffer_0_37 : _GEN_1831; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1833 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_5_T_3[5:0] ? buffer_0_38 : _GEN_1832; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1834 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_5_T_3[5:0] ? buffer_0_39 : _GEN_1833; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1835 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_5_T_3[5:0] ? buffer_0_40 : _GEN_1834; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1836 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_5_T_3[5:0] ? buffer_0_41 : _GEN_1835; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1837 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_5_T_3[5:0] ? buffer_0_42 : _GEN_1836; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1838 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_5_T_3[5:0] ? buffer_0_43 : _GEN_1837; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1839 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_5_T_3[5:0] ? buffer_0_44 : _GEN_1838; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1840 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_5_T_3[5:0] ? buffer_0_45 : _GEN_1839; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1841 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_5_T_3[5:0] ? buffer_0_46 : _GEN_1840; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1842 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_5_T_3[5:0] ? buffer_0_47 : _GEN_1841; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1843 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_5_T_3[5:0] ? buffer_0_48 : _GEN_1842; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1844 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_5_T_3[5:0] ? buffer_0_49 : _GEN_1843; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1845 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_5_T_3[5:0] ? buffer_0_50 : _GEN_1844; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1846 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_5_T_3[5:0] ? buffer_0_51 : _GEN_1845; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1847 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_5_T_3[5:0] ? buffer_0_52 : _GEN_1846; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1848 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_5_T_3[5:0] ? buffer_0_53 : _GEN_1847; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1849 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_5_T_3[5:0] ? buffer_0_54 : _GEN_1848; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1850 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_5_T_3[5:0] ? buffer_0_55 : _GEN_1849; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1851 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_5_T_3[5:0] ? buffer_0_56 : _GEN_1850; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1852 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_5_T_3[5:0] ? buffer_0_57 : _GEN_1851; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1853 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_5_T_3[5:0] ? buffer_0_58 : _GEN_1852; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1854 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_5_T_3[5:0] ? buffer_0_59 : _GEN_1853; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1855 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_5_T_3[5:0] ? buffer_0_60 : _GEN_1854; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1856 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_5_T_3[5:0] ? buffer_0_61 : _GEN_1855; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1857 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_5_T_3[5:0] ? buffer_0_62 : _GEN_1856; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1858 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_5_T_3[5:0] ? buffer_0_63 : _GEN_1857; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1859 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_5_T_3[5:0] ? buffer_1_0 : _GEN_1858; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1860 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_5_T_3[5:0] ? buffer_1_1 : _GEN_1859; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1861 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_5_T_3[5:0] ? buffer_1_2 : _GEN_1860; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1862 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_5_T_3[5:0] ? buffer_1_3 : _GEN_1861; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1863 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_5_T_3[5:0] ? buffer_1_4 : _GEN_1862; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1864 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_5_T_3[5:0] ? buffer_1_5 : _GEN_1863; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1865 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_5_T_3[5:0] ? buffer_1_6 : _GEN_1864; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1866 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_5_T_3[5:0] ? buffer_1_7 : _GEN_1865; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1867 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_5_T_3[5:0] ? buffer_1_8 : _GEN_1866; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1868 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_5_T_3[5:0] ? buffer_1_9 : _GEN_1867; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1869 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_5_T_3[5:0] ? buffer_1_10 : _GEN_1868; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1870 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_5_T_3[5:0] ? buffer_1_11 : _GEN_1869; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1871 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_5_T_3[5:0] ? buffer_1_12 : _GEN_1870; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1872 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_5_T_3[5:0] ? buffer_1_13 : _GEN_1871; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1873 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_5_T_3[5:0] ? buffer_1_14 : _GEN_1872; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1874 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_5_T_3[5:0] ? buffer_1_15 : _GEN_1873; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1875 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_5_T_3[5:0] ? buffer_1_16 : _GEN_1874; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1876 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_5_T_3[5:0] ? buffer_1_17 : _GEN_1875; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1877 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_5_T_3[5:0] ? buffer_1_18 : _GEN_1876; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1878 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_5_T_3[5:0] ? buffer_1_19 : _GEN_1877; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1879 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_5_T_3[5:0] ? buffer_1_20 : _GEN_1878; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1880 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_5_T_3[5:0] ? buffer_1_21 : _GEN_1879; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1881 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_5_T_3[5:0] ? buffer_1_22 : _GEN_1880; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1882 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_5_T_3[5:0] ? buffer_1_23 : _GEN_1881; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1883 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_5_T_3[5:0] ? buffer_1_24 : _GEN_1882; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1884 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_5_T_3[5:0] ? buffer_1_25 : _GEN_1883; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1885 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_5_T_3[5:0] ? buffer_1_26 : _GEN_1884; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1886 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_5_T_3[5:0] ? buffer_1_27 : _GEN_1885; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1887 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_5_T_3[5:0] ? buffer_1_28 : _GEN_1886; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1888 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_5_T_3[5:0] ? buffer_1_29 : _GEN_1887; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1889 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_5_T_3[5:0] ? buffer_1_30 : _GEN_1888; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1890 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_5_T_3[5:0] ? buffer_1_31 : _GEN_1889; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1891 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_5_T_3[5:0] ? buffer_1_32 : _GEN_1890; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1892 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_5_T_3[5:0] ? buffer_1_33 : _GEN_1891; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1893 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_5_T_3[5:0] ? buffer_1_34 : _GEN_1892; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1894 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_5_T_3[5:0] ? buffer_1_35 : _GEN_1893; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1895 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_5_T_3[5:0] ? buffer_1_36 : _GEN_1894; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1896 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_5_T_3[5:0] ? buffer_1_37 : _GEN_1895; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1897 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_5_T_3[5:0] ? buffer_1_38 : _GEN_1896; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1898 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_5_T_3[5:0] ? buffer_1_39 : _GEN_1897; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1899 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_5_T_3[5:0] ? buffer_1_40 : _GEN_1898; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1900 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_5_T_3[5:0] ? buffer_1_41 : _GEN_1899; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1901 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_5_T_3[5:0] ? buffer_1_42 : _GEN_1900; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1902 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_5_T_3[5:0] ? buffer_1_43 : _GEN_1901; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1903 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_5_T_3[5:0] ? buffer_1_44 : _GEN_1902; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1904 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_5_T_3[5:0] ? buffer_1_45 : _GEN_1903; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1905 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_5_T_3[5:0] ? buffer_1_46 : _GEN_1904; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1906 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_5_T_3[5:0] ? buffer_1_47 : _GEN_1905; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1907 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_5_T_3[5:0] ? buffer_1_48 : _GEN_1906; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1908 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_5_T_3[5:0] ? buffer_1_49 : _GEN_1907; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1909 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_5_T_3[5:0] ? buffer_1_50 : _GEN_1908; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1910 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_5_T_3[5:0] ? buffer_1_51 : _GEN_1909; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1911 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_5_T_3[5:0] ? buffer_1_52 : _GEN_1910; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1912 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_5_T_3[5:0] ? buffer_1_53 : _GEN_1911; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1913 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_5_T_3[5:0] ? buffer_1_54 : _GEN_1912; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1914 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_5_T_3[5:0] ? buffer_1_55 : _GEN_1913; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1915 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_5_T_3[5:0] ? buffer_1_56 : _GEN_1914; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1916 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_5_T_3[5:0] ? buffer_1_57 : _GEN_1915; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1917 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_5_T_3[5:0] ? buffer_1_58 : _GEN_1916; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1918 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_5_T_3[5:0] ? buffer_1_59 : _GEN_1917; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1919 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_5_T_3[5:0] ? buffer_1_60 : _GEN_1918; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1920 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_5_T_3[5:0] ? buffer_1_61 : _GEN_1919; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1921 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_5_T_3[5:0] ? buffer_1_62 : _GEN_1920; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1922 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_5_T_3[5:0] ? buffer_1_63 : _GEN_1921; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1923 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_5_T_3[5:0] ? buffer_2_0 : _GEN_1922; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1924 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_5_T_3[5:0] ? buffer_2_1 : _GEN_1923; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1925 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_5_T_3[5:0] ? buffer_2_2 : _GEN_1924; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1926 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_5_T_3[5:0] ? buffer_2_3 : _GEN_1925; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1927 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_5_T_3[5:0] ? buffer_2_4 : _GEN_1926; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1928 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_5_T_3[5:0] ? buffer_2_5 : _GEN_1927; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1929 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_5_T_3[5:0] ? buffer_2_6 : _GEN_1928; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1930 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_5_T_3[5:0] ? buffer_2_7 : _GEN_1929; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1931 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_5_T_3[5:0] ? buffer_2_8 : _GEN_1930; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1932 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_5_T_3[5:0] ? buffer_2_9 : _GEN_1931; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1933 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_5_T_3[5:0] ? buffer_2_10 : _GEN_1932; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1934 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_5_T_3[5:0] ? buffer_2_11 : _GEN_1933; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1935 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_5_T_3[5:0] ? buffer_2_12 : _GEN_1934; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1936 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_5_T_3[5:0] ? buffer_2_13 : _GEN_1935; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1937 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_5_T_3[5:0] ? buffer_2_14 : _GEN_1936; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1938 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_5_T_3[5:0] ? buffer_2_15 : _GEN_1937; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1939 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_5_T_3[5:0] ? buffer_2_16 : _GEN_1938; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1940 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_5_T_3[5:0] ? buffer_2_17 : _GEN_1939; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1941 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_5_T_3[5:0] ? buffer_2_18 : _GEN_1940; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1942 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_5_T_3[5:0] ? buffer_2_19 : _GEN_1941; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1943 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_5_T_3[5:0] ? buffer_2_20 : _GEN_1942; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1944 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_5_T_3[5:0] ? buffer_2_21 : _GEN_1943; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1945 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_5_T_3[5:0] ? buffer_2_22 : _GEN_1944; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1946 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_5_T_3[5:0] ? buffer_2_23 : _GEN_1945; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1947 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_5_T_3[5:0] ? buffer_2_24 : _GEN_1946; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1948 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_5_T_3[5:0] ? buffer_2_25 : _GEN_1947; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1949 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_5_T_3[5:0] ? buffer_2_26 : _GEN_1948; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1950 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_5_T_3[5:0] ? buffer_2_27 : _GEN_1949; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1951 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_5_T_3[5:0] ? buffer_2_28 : _GEN_1950; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1952 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_5_T_3[5:0] ? buffer_2_29 : _GEN_1951; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1953 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_5_T_3[5:0] ? buffer_2_30 : _GEN_1952; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1954 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_5_T_3[5:0] ? buffer_2_31 : _GEN_1953; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1955 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_5_T_3[5:0] ? buffer_2_32 : _GEN_1954; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1956 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_5_T_3[5:0] ? buffer_2_33 : _GEN_1955; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1957 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_5_T_3[5:0] ? buffer_2_34 : _GEN_1956; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1958 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_5_T_3[5:0] ? buffer_2_35 : _GEN_1957; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1959 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_5_T_3[5:0] ? buffer_2_36 : _GEN_1958; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1960 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_5_T_3[5:0] ? buffer_2_37 : _GEN_1959; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1961 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_5_T_3[5:0] ? buffer_2_38 : _GEN_1960; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1962 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_5_T_3[5:0] ? buffer_2_39 : _GEN_1961; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1963 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_5_T_3[5:0] ? buffer_2_40 : _GEN_1962; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1964 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_5_T_3[5:0] ? buffer_2_41 : _GEN_1963; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1965 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_5_T_3[5:0] ? buffer_2_42 : _GEN_1964; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1966 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_5_T_3[5:0] ? buffer_2_43 : _GEN_1965; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1967 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_5_T_3[5:0] ? buffer_2_44 : _GEN_1966; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1968 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_5_T_3[5:0] ? buffer_2_45 : _GEN_1967; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1969 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_5_T_3[5:0] ? buffer_2_46 : _GEN_1968; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1970 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_5_T_3[5:0] ? buffer_2_47 : _GEN_1969; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1971 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_5_T_3[5:0] ? buffer_2_48 : _GEN_1970; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1972 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_5_T_3[5:0] ? buffer_2_49 : _GEN_1971; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1973 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_5_T_3[5:0] ? buffer_2_50 : _GEN_1972; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1974 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_5_T_3[5:0] ? buffer_2_51 : _GEN_1973; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1975 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_5_T_3[5:0] ? buffer_2_52 : _GEN_1974; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1976 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_5_T_3[5:0] ? buffer_2_53 : _GEN_1975; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1977 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_5_T_3[5:0] ? buffer_2_54 : _GEN_1976; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1978 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_5_T_3[5:0] ? buffer_2_55 : _GEN_1977; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1979 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_5_T_3[5:0] ? buffer_2_56 : _GEN_1978; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1980 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_5_T_3[5:0] ? buffer_2_57 : _GEN_1979; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1981 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_5_T_3[5:0] ? buffer_2_58 : _GEN_1980; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1982 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_5_T_3[5:0] ? buffer_2_59 : _GEN_1981; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1983 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_5_T_3[5:0] ? buffer_2_60 : _GEN_1982; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1984 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_5_T_3[5:0] ? buffer_2_61 : _GEN_1983; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1985 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_5_T_3[5:0] ? buffer_2_62 : _GEN_1984; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1986 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_5_T_3[5:0] ? buffer_2_63 : _GEN_1985; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1987 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_5_T_3[5:0] ? buffer_3_0 : _GEN_1986; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1988 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_5_T_3[5:0] ? buffer_3_1 : _GEN_1987; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1989 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_5_T_3[5:0] ? buffer_3_2 : _GEN_1988; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1990 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_5_T_3[5:0] ? buffer_3_3 : _GEN_1989; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1991 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_5_T_3[5:0] ? buffer_3_4 : _GEN_1990; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1992 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_5_T_3[5:0] ? buffer_3_5 : _GEN_1991; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1993 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_5_T_3[5:0] ? buffer_3_6 : _GEN_1992; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1994 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_5_T_3[5:0] ? buffer_3_7 : _GEN_1993; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1995 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_5_T_3[5:0] ? buffer_3_8 : _GEN_1994; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1996 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_5_T_3[5:0] ? buffer_3_9 : _GEN_1995; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1997 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_5_T_3[5:0] ? buffer_3_10 : _GEN_1996; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1998 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_5_T_3[5:0] ? buffer_3_11 : _GEN_1997; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_1999 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_5_T_3[5:0] ? buffer_3_12 : _GEN_1998; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2000 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_5_T_3[5:0] ? buffer_3_13 : _GEN_1999; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2001 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_5_T_3[5:0] ? buffer_3_14 : _GEN_2000; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2002 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_5_T_3[5:0] ? buffer_3_15 : _GEN_2001; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2003 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_5_T_3[5:0] ? buffer_3_16 : _GEN_2002; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2004 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_5_T_3[5:0] ? buffer_3_17 : _GEN_2003; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2005 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_5_T_3[5:0] ? buffer_3_18 : _GEN_2004; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2006 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_5_T_3[5:0] ? buffer_3_19 : _GEN_2005; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2007 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_5_T_3[5:0] ? buffer_3_20 : _GEN_2006; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2008 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_5_T_3[5:0] ? buffer_3_21 : _GEN_2007; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2009 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_5_T_3[5:0] ? buffer_3_22 : _GEN_2008; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2010 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_5_T_3[5:0] ? buffer_3_23 : _GEN_2009; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2011 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_5_T_3[5:0] ? buffer_3_24 : _GEN_2010; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2012 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_5_T_3[5:0] ? buffer_3_25 : _GEN_2011; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2013 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_5_T_3[5:0] ? buffer_3_26 : _GEN_2012; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2014 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_5_T_3[5:0] ? buffer_3_27 : _GEN_2013; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2015 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_5_T_3[5:0] ? buffer_3_28 : _GEN_2014; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2016 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_5_T_3[5:0] ? buffer_3_29 : _GEN_2015; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2017 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_5_T_3[5:0] ? buffer_3_30 : _GEN_2016; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2018 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_5_T_3[5:0] ? buffer_3_31 : _GEN_2017; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2019 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_5_T_3[5:0] ? buffer_3_32 : _GEN_2018; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2020 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_5_T_3[5:0] ? buffer_3_33 : _GEN_2019; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2021 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_5_T_3[5:0] ? buffer_3_34 : _GEN_2020; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2022 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_5_T_3[5:0] ? buffer_3_35 : _GEN_2021; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2023 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_5_T_3[5:0] ? buffer_3_36 : _GEN_2022; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2024 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_5_T_3[5:0] ? buffer_3_37 : _GEN_2023; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2025 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_5_T_3[5:0] ? buffer_3_38 : _GEN_2024; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2026 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_5_T_3[5:0] ? buffer_3_39 : _GEN_2025; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2027 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_5_T_3[5:0] ? buffer_3_40 : _GEN_2026; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2028 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_5_T_3[5:0] ? buffer_3_41 : _GEN_2027; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2029 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_5_T_3[5:0] ? buffer_3_42 : _GEN_2028; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2030 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_5_T_3[5:0] ? buffer_3_43 : _GEN_2029; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2031 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_5_T_3[5:0] ? buffer_3_44 : _GEN_2030; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2032 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_5_T_3[5:0] ? buffer_3_45 : _GEN_2031; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2033 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_5_T_3[5:0] ? buffer_3_46 : _GEN_2032; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2034 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_5_T_3[5:0] ? buffer_3_47 : _GEN_2033; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2035 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_5_T_3[5:0] ? buffer_3_48 : _GEN_2034; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2036 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_5_T_3[5:0] ? buffer_3_49 : _GEN_2035; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2037 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_5_T_3[5:0] ? buffer_3_50 : _GEN_2036; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2038 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_5_T_3[5:0] ? buffer_3_51 : _GEN_2037; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2039 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_5_T_3[5:0] ? buffer_3_52 : _GEN_2038; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2040 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_5_T_3[5:0] ? buffer_3_53 : _GEN_2039; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2041 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_5_T_3[5:0] ? buffer_3_54 : _GEN_2040; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2042 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_5_T_3[5:0] ? buffer_3_55 : _GEN_2041; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2043 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_5_T_3[5:0] ? buffer_3_56 : _GEN_2042; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2044 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_5_T_3[5:0] ? buffer_3_57 : _GEN_2043; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2045 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_5_T_3[5:0] ? buffer_3_58 : _GEN_2044; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2046 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_5_T_3[5:0] ? buffer_3_59 : _GEN_2045; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2047 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_5_T_3[5:0] ? buffer_3_60 : _GEN_2046; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2048 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_5_T_3[5:0] ? buffer_3_61 : _GEN_2047; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2049 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_5_T_3[5:0] ? buffer_3_62 : _GEN_2048; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2050 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_5_T_3[5:0] ? buffer_3_63 : _GEN_2049; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_6_T_3 = _io_out_weight_0_T_1 + 8'h6; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_2052 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_6_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2053 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_6_T_3[5:0] ? buffer_0_2 : _GEN_2052; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2054 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_6_T_3[5:0] ? buffer_0_3 : _GEN_2053; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2055 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_6_T_3[5:0] ? buffer_0_4 : _GEN_2054; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2056 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_6_T_3[5:0] ? buffer_0_5 : _GEN_2055; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2057 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_6_T_3[5:0] ? buffer_0_6 : _GEN_2056; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2058 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_6_T_3[5:0] ? buffer_0_7 : _GEN_2057; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2059 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_6_T_3[5:0] ? buffer_0_8 : _GEN_2058; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2060 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_6_T_3[5:0] ? buffer_0_9 : _GEN_2059; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2061 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_6_T_3[5:0] ? buffer_0_10 : _GEN_2060; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2062 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_6_T_3[5:0] ? buffer_0_11 : _GEN_2061; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2063 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_6_T_3[5:0] ? buffer_0_12 : _GEN_2062; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2064 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_6_T_3[5:0] ? buffer_0_13 : _GEN_2063; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2065 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_6_T_3[5:0] ? buffer_0_14 : _GEN_2064; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2066 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_6_T_3[5:0] ? buffer_0_15 : _GEN_2065; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2067 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_6_T_3[5:0] ? buffer_0_16 : _GEN_2066; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2068 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_6_T_3[5:0] ? buffer_0_17 : _GEN_2067; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2069 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_6_T_3[5:0] ? buffer_0_18 : _GEN_2068; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2070 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_6_T_3[5:0] ? buffer_0_19 : _GEN_2069; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2071 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_6_T_3[5:0] ? buffer_0_20 : _GEN_2070; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2072 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_6_T_3[5:0] ? buffer_0_21 : _GEN_2071; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2073 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_6_T_3[5:0] ? buffer_0_22 : _GEN_2072; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2074 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_6_T_3[5:0] ? buffer_0_23 : _GEN_2073; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2075 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_6_T_3[5:0] ? buffer_0_24 : _GEN_2074; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2076 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_6_T_3[5:0] ? buffer_0_25 : _GEN_2075; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2077 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_6_T_3[5:0] ? buffer_0_26 : _GEN_2076; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2078 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_6_T_3[5:0] ? buffer_0_27 : _GEN_2077; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2079 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_6_T_3[5:0] ? buffer_0_28 : _GEN_2078; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2080 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_6_T_3[5:0] ? buffer_0_29 : _GEN_2079; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2081 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_6_T_3[5:0] ? buffer_0_30 : _GEN_2080; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2082 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_6_T_3[5:0] ? buffer_0_31 : _GEN_2081; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2083 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_6_T_3[5:0] ? buffer_0_32 : _GEN_2082; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2084 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_6_T_3[5:0] ? buffer_0_33 : _GEN_2083; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2085 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_6_T_3[5:0] ? buffer_0_34 : _GEN_2084; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2086 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_6_T_3[5:0] ? buffer_0_35 : _GEN_2085; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2087 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_6_T_3[5:0] ? buffer_0_36 : _GEN_2086; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2088 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_6_T_3[5:0] ? buffer_0_37 : _GEN_2087; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2089 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_6_T_3[5:0] ? buffer_0_38 : _GEN_2088; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2090 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_6_T_3[5:0] ? buffer_0_39 : _GEN_2089; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2091 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_6_T_3[5:0] ? buffer_0_40 : _GEN_2090; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2092 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_6_T_3[5:0] ? buffer_0_41 : _GEN_2091; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2093 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_6_T_3[5:0] ? buffer_0_42 : _GEN_2092; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2094 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_6_T_3[5:0] ? buffer_0_43 : _GEN_2093; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2095 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_6_T_3[5:0] ? buffer_0_44 : _GEN_2094; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2096 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_6_T_3[5:0] ? buffer_0_45 : _GEN_2095; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2097 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_6_T_3[5:0] ? buffer_0_46 : _GEN_2096; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2098 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_6_T_3[5:0] ? buffer_0_47 : _GEN_2097; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2099 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_6_T_3[5:0] ? buffer_0_48 : _GEN_2098; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2100 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_6_T_3[5:0] ? buffer_0_49 : _GEN_2099; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2101 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_6_T_3[5:0] ? buffer_0_50 : _GEN_2100; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2102 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_6_T_3[5:0] ? buffer_0_51 : _GEN_2101; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2103 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_6_T_3[5:0] ? buffer_0_52 : _GEN_2102; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2104 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_6_T_3[5:0] ? buffer_0_53 : _GEN_2103; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2105 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_6_T_3[5:0] ? buffer_0_54 : _GEN_2104; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2106 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_6_T_3[5:0] ? buffer_0_55 : _GEN_2105; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2107 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_6_T_3[5:0] ? buffer_0_56 : _GEN_2106; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2108 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_6_T_3[5:0] ? buffer_0_57 : _GEN_2107; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2109 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_6_T_3[5:0] ? buffer_0_58 : _GEN_2108; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2110 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_6_T_3[5:0] ? buffer_0_59 : _GEN_2109; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2111 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_6_T_3[5:0] ? buffer_0_60 : _GEN_2110; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2112 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_6_T_3[5:0] ? buffer_0_61 : _GEN_2111; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2113 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_6_T_3[5:0] ? buffer_0_62 : _GEN_2112; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2114 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_6_T_3[5:0] ? buffer_0_63 : _GEN_2113; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2115 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_6_T_3[5:0] ? buffer_1_0 : _GEN_2114; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2116 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_6_T_3[5:0] ? buffer_1_1 : _GEN_2115; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2117 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_6_T_3[5:0] ? buffer_1_2 : _GEN_2116; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2118 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_6_T_3[5:0] ? buffer_1_3 : _GEN_2117; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2119 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_6_T_3[5:0] ? buffer_1_4 : _GEN_2118; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2120 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_6_T_3[5:0] ? buffer_1_5 : _GEN_2119; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2121 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_6_T_3[5:0] ? buffer_1_6 : _GEN_2120; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2122 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_6_T_3[5:0] ? buffer_1_7 : _GEN_2121; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2123 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_6_T_3[5:0] ? buffer_1_8 : _GEN_2122; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2124 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_6_T_3[5:0] ? buffer_1_9 : _GEN_2123; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2125 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_6_T_3[5:0] ? buffer_1_10 : _GEN_2124; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2126 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_6_T_3[5:0] ? buffer_1_11 : _GEN_2125; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2127 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_6_T_3[5:0] ? buffer_1_12 : _GEN_2126; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2128 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_6_T_3[5:0] ? buffer_1_13 : _GEN_2127; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2129 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_6_T_3[5:0] ? buffer_1_14 : _GEN_2128; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2130 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_6_T_3[5:0] ? buffer_1_15 : _GEN_2129; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2131 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_6_T_3[5:0] ? buffer_1_16 : _GEN_2130; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2132 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_6_T_3[5:0] ? buffer_1_17 : _GEN_2131; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2133 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_6_T_3[5:0] ? buffer_1_18 : _GEN_2132; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2134 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_6_T_3[5:0] ? buffer_1_19 : _GEN_2133; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2135 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_6_T_3[5:0] ? buffer_1_20 : _GEN_2134; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2136 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_6_T_3[5:0] ? buffer_1_21 : _GEN_2135; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2137 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_6_T_3[5:0] ? buffer_1_22 : _GEN_2136; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2138 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_6_T_3[5:0] ? buffer_1_23 : _GEN_2137; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2139 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_6_T_3[5:0] ? buffer_1_24 : _GEN_2138; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2140 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_6_T_3[5:0] ? buffer_1_25 : _GEN_2139; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2141 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_6_T_3[5:0] ? buffer_1_26 : _GEN_2140; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2142 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_6_T_3[5:0] ? buffer_1_27 : _GEN_2141; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2143 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_6_T_3[5:0] ? buffer_1_28 : _GEN_2142; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2144 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_6_T_3[5:0] ? buffer_1_29 : _GEN_2143; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2145 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_6_T_3[5:0] ? buffer_1_30 : _GEN_2144; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2146 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_6_T_3[5:0] ? buffer_1_31 : _GEN_2145; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2147 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_6_T_3[5:0] ? buffer_1_32 : _GEN_2146; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2148 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_6_T_3[5:0] ? buffer_1_33 : _GEN_2147; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2149 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_6_T_3[5:0] ? buffer_1_34 : _GEN_2148; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2150 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_6_T_3[5:0] ? buffer_1_35 : _GEN_2149; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2151 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_6_T_3[5:0] ? buffer_1_36 : _GEN_2150; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2152 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_6_T_3[5:0] ? buffer_1_37 : _GEN_2151; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2153 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_6_T_3[5:0] ? buffer_1_38 : _GEN_2152; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2154 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_6_T_3[5:0] ? buffer_1_39 : _GEN_2153; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2155 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_6_T_3[5:0] ? buffer_1_40 : _GEN_2154; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2156 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_6_T_3[5:0] ? buffer_1_41 : _GEN_2155; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2157 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_6_T_3[5:0] ? buffer_1_42 : _GEN_2156; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2158 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_6_T_3[5:0] ? buffer_1_43 : _GEN_2157; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2159 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_6_T_3[5:0] ? buffer_1_44 : _GEN_2158; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2160 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_6_T_3[5:0] ? buffer_1_45 : _GEN_2159; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2161 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_6_T_3[5:0] ? buffer_1_46 : _GEN_2160; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2162 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_6_T_3[5:0] ? buffer_1_47 : _GEN_2161; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2163 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_6_T_3[5:0] ? buffer_1_48 : _GEN_2162; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2164 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_6_T_3[5:0] ? buffer_1_49 : _GEN_2163; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2165 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_6_T_3[5:0] ? buffer_1_50 : _GEN_2164; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2166 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_6_T_3[5:0] ? buffer_1_51 : _GEN_2165; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2167 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_6_T_3[5:0] ? buffer_1_52 : _GEN_2166; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2168 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_6_T_3[5:0] ? buffer_1_53 : _GEN_2167; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2169 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_6_T_3[5:0] ? buffer_1_54 : _GEN_2168; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2170 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_6_T_3[5:0] ? buffer_1_55 : _GEN_2169; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2171 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_6_T_3[5:0] ? buffer_1_56 : _GEN_2170; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2172 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_6_T_3[5:0] ? buffer_1_57 : _GEN_2171; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2173 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_6_T_3[5:0] ? buffer_1_58 : _GEN_2172; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2174 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_6_T_3[5:0] ? buffer_1_59 : _GEN_2173; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2175 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_6_T_3[5:0] ? buffer_1_60 : _GEN_2174; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2176 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_6_T_3[5:0] ? buffer_1_61 : _GEN_2175; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2177 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_6_T_3[5:0] ? buffer_1_62 : _GEN_2176; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2178 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_6_T_3[5:0] ? buffer_1_63 : _GEN_2177; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2179 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_6_T_3[5:0] ? buffer_2_0 : _GEN_2178; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2180 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_6_T_3[5:0] ? buffer_2_1 : _GEN_2179; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2181 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_6_T_3[5:0] ? buffer_2_2 : _GEN_2180; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2182 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_6_T_3[5:0] ? buffer_2_3 : _GEN_2181; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2183 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_6_T_3[5:0] ? buffer_2_4 : _GEN_2182; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2184 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_6_T_3[5:0] ? buffer_2_5 : _GEN_2183; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2185 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_6_T_3[5:0] ? buffer_2_6 : _GEN_2184; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2186 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_6_T_3[5:0] ? buffer_2_7 : _GEN_2185; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2187 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_6_T_3[5:0] ? buffer_2_8 : _GEN_2186; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2188 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_6_T_3[5:0] ? buffer_2_9 : _GEN_2187; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2189 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_6_T_3[5:0] ? buffer_2_10 : _GEN_2188; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2190 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_6_T_3[5:0] ? buffer_2_11 : _GEN_2189; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2191 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_6_T_3[5:0] ? buffer_2_12 : _GEN_2190; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2192 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_6_T_3[5:0] ? buffer_2_13 : _GEN_2191; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2193 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_6_T_3[5:0] ? buffer_2_14 : _GEN_2192; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2194 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_6_T_3[5:0] ? buffer_2_15 : _GEN_2193; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2195 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_6_T_3[5:0] ? buffer_2_16 : _GEN_2194; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2196 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_6_T_3[5:0] ? buffer_2_17 : _GEN_2195; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2197 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_6_T_3[5:0] ? buffer_2_18 : _GEN_2196; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2198 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_6_T_3[5:0] ? buffer_2_19 : _GEN_2197; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2199 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_6_T_3[5:0] ? buffer_2_20 : _GEN_2198; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2200 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_6_T_3[5:0] ? buffer_2_21 : _GEN_2199; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2201 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_6_T_3[5:0] ? buffer_2_22 : _GEN_2200; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2202 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_6_T_3[5:0] ? buffer_2_23 : _GEN_2201; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2203 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_6_T_3[5:0] ? buffer_2_24 : _GEN_2202; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2204 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_6_T_3[5:0] ? buffer_2_25 : _GEN_2203; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2205 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_6_T_3[5:0] ? buffer_2_26 : _GEN_2204; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2206 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_6_T_3[5:0] ? buffer_2_27 : _GEN_2205; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2207 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_6_T_3[5:0] ? buffer_2_28 : _GEN_2206; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2208 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_6_T_3[5:0] ? buffer_2_29 : _GEN_2207; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2209 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_6_T_3[5:0] ? buffer_2_30 : _GEN_2208; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2210 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_6_T_3[5:0] ? buffer_2_31 : _GEN_2209; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2211 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_6_T_3[5:0] ? buffer_2_32 : _GEN_2210; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2212 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_6_T_3[5:0] ? buffer_2_33 : _GEN_2211; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2213 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_6_T_3[5:0] ? buffer_2_34 : _GEN_2212; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2214 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_6_T_3[5:0] ? buffer_2_35 : _GEN_2213; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2215 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_6_T_3[5:0] ? buffer_2_36 : _GEN_2214; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2216 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_6_T_3[5:0] ? buffer_2_37 : _GEN_2215; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2217 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_6_T_3[5:0] ? buffer_2_38 : _GEN_2216; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2218 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_6_T_3[5:0] ? buffer_2_39 : _GEN_2217; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2219 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_6_T_3[5:0] ? buffer_2_40 : _GEN_2218; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2220 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_6_T_3[5:0] ? buffer_2_41 : _GEN_2219; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2221 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_6_T_3[5:0] ? buffer_2_42 : _GEN_2220; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2222 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_6_T_3[5:0] ? buffer_2_43 : _GEN_2221; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2223 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_6_T_3[5:0] ? buffer_2_44 : _GEN_2222; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2224 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_6_T_3[5:0] ? buffer_2_45 : _GEN_2223; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2225 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_6_T_3[5:0] ? buffer_2_46 : _GEN_2224; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2226 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_6_T_3[5:0] ? buffer_2_47 : _GEN_2225; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2227 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_6_T_3[5:0] ? buffer_2_48 : _GEN_2226; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2228 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_6_T_3[5:0] ? buffer_2_49 : _GEN_2227; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2229 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_6_T_3[5:0] ? buffer_2_50 : _GEN_2228; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2230 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_6_T_3[5:0] ? buffer_2_51 : _GEN_2229; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2231 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_6_T_3[5:0] ? buffer_2_52 : _GEN_2230; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2232 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_6_T_3[5:0] ? buffer_2_53 : _GEN_2231; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2233 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_6_T_3[5:0] ? buffer_2_54 : _GEN_2232; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2234 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_6_T_3[5:0] ? buffer_2_55 : _GEN_2233; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2235 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_6_T_3[5:0] ? buffer_2_56 : _GEN_2234; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2236 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_6_T_3[5:0] ? buffer_2_57 : _GEN_2235; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2237 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_6_T_3[5:0] ? buffer_2_58 : _GEN_2236; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2238 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_6_T_3[5:0] ? buffer_2_59 : _GEN_2237; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2239 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_6_T_3[5:0] ? buffer_2_60 : _GEN_2238; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2240 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_6_T_3[5:0] ? buffer_2_61 : _GEN_2239; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2241 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_6_T_3[5:0] ? buffer_2_62 : _GEN_2240; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2242 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_6_T_3[5:0] ? buffer_2_63 : _GEN_2241; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2243 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_6_T_3[5:0] ? buffer_3_0 : _GEN_2242; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2244 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_6_T_3[5:0] ? buffer_3_1 : _GEN_2243; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2245 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_6_T_3[5:0] ? buffer_3_2 : _GEN_2244; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2246 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_6_T_3[5:0] ? buffer_3_3 : _GEN_2245; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2247 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_6_T_3[5:0] ? buffer_3_4 : _GEN_2246; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2248 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_6_T_3[5:0] ? buffer_3_5 : _GEN_2247; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2249 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_6_T_3[5:0] ? buffer_3_6 : _GEN_2248; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2250 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_6_T_3[5:0] ? buffer_3_7 : _GEN_2249; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2251 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_6_T_3[5:0] ? buffer_3_8 : _GEN_2250; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2252 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_6_T_3[5:0] ? buffer_3_9 : _GEN_2251; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2253 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_6_T_3[5:0] ? buffer_3_10 : _GEN_2252; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2254 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_6_T_3[5:0] ? buffer_3_11 : _GEN_2253; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2255 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_6_T_3[5:0] ? buffer_3_12 : _GEN_2254; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2256 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_6_T_3[5:0] ? buffer_3_13 : _GEN_2255; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2257 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_6_T_3[5:0] ? buffer_3_14 : _GEN_2256; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2258 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_6_T_3[5:0] ? buffer_3_15 : _GEN_2257; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2259 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_6_T_3[5:0] ? buffer_3_16 : _GEN_2258; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2260 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_6_T_3[5:0] ? buffer_3_17 : _GEN_2259; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2261 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_6_T_3[5:0] ? buffer_3_18 : _GEN_2260; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2262 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_6_T_3[5:0] ? buffer_3_19 : _GEN_2261; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2263 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_6_T_3[5:0] ? buffer_3_20 : _GEN_2262; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2264 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_6_T_3[5:0] ? buffer_3_21 : _GEN_2263; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2265 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_6_T_3[5:0] ? buffer_3_22 : _GEN_2264; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2266 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_6_T_3[5:0] ? buffer_3_23 : _GEN_2265; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2267 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_6_T_3[5:0] ? buffer_3_24 : _GEN_2266; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2268 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_6_T_3[5:0] ? buffer_3_25 : _GEN_2267; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2269 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_6_T_3[5:0] ? buffer_3_26 : _GEN_2268; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2270 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_6_T_3[5:0] ? buffer_3_27 : _GEN_2269; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2271 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_6_T_3[5:0] ? buffer_3_28 : _GEN_2270; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2272 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_6_T_3[5:0] ? buffer_3_29 : _GEN_2271; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2273 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_6_T_3[5:0] ? buffer_3_30 : _GEN_2272; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2274 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_6_T_3[5:0] ? buffer_3_31 : _GEN_2273; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2275 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_6_T_3[5:0] ? buffer_3_32 : _GEN_2274; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2276 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_6_T_3[5:0] ? buffer_3_33 : _GEN_2275; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2277 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_6_T_3[5:0] ? buffer_3_34 : _GEN_2276; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2278 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_6_T_3[5:0] ? buffer_3_35 : _GEN_2277; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2279 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_6_T_3[5:0] ? buffer_3_36 : _GEN_2278; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2280 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_6_T_3[5:0] ? buffer_3_37 : _GEN_2279; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2281 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_6_T_3[5:0] ? buffer_3_38 : _GEN_2280; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2282 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_6_T_3[5:0] ? buffer_3_39 : _GEN_2281; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2283 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_6_T_3[5:0] ? buffer_3_40 : _GEN_2282; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2284 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_6_T_3[5:0] ? buffer_3_41 : _GEN_2283; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2285 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_6_T_3[5:0] ? buffer_3_42 : _GEN_2284; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2286 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_6_T_3[5:0] ? buffer_3_43 : _GEN_2285; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2287 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_6_T_3[5:0] ? buffer_3_44 : _GEN_2286; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2288 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_6_T_3[5:0] ? buffer_3_45 : _GEN_2287; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2289 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_6_T_3[5:0] ? buffer_3_46 : _GEN_2288; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2290 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_6_T_3[5:0] ? buffer_3_47 : _GEN_2289; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2291 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_6_T_3[5:0] ? buffer_3_48 : _GEN_2290; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2292 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_6_T_3[5:0] ? buffer_3_49 : _GEN_2291; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2293 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_6_T_3[5:0] ? buffer_3_50 : _GEN_2292; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2294 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_6_T_3[5:0] ? buffer_3_51 : _GEN_2293; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2295 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_6_T_3[5:0] ? buffer_3_52 : _GEN_2294; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2296 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_6_T_3[5:0] ? buffer_3_53 : _GEN_2295; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2297 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_6_T_3[5:0] ? buffer_3_54 : _GEN_2296; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2298 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_6_T_3[5:0] ? buffer_3_55 : _GEN_2297; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2299 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_6_T_3[5:0] ? buffer_3_56 : _GEN_2298; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2300 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_6_T_3[5:0] ? buffer_3_57 : _GEN_2299; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2301 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_6_T_3[5:0] ? buffer_3_58 : _GEN_2300; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2302 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_6_T_3[5:0] ? buffer_3_59 : _GEN_2301; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2303 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_6_T_3[5:0] ? buffer_3_60 : _GEN_2302; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2304 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_6_T_3[5:0] ? buffer_3_61 : _GEN_2303; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2305 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_6_T_3[5:0] ? buffer_3_62 : _GEN_2304; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2306 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_6_T_3[5:0] ? buffer_3_63 : _GEN_2305; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _io_out_weight_7_T_3 = _io_out_weight_0_T_1 + 8'h7; // @[Weight_Buffer.scala 64:88]
  wire [7:0] _GEN_2308 = 2'h0 == read_ptr[1:0] & 6'h1 == _io_out_weight_7_T_3[5:0] ? buffer_0_1 : buffer_0_0; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2309 = 2'h0 == read_ptr[1:0] & 6'h2 == _io_out_weight_7_T_3[5:0] ? buffer_0_2 : _GEN_2308; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2310 = 2'h0 == read_ptr[1:0] & 6'h3 == _io_out_weight_7_T_3[5:0] ? buffer_0_3 : _GEN_2309; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2311 = 2'h0 == read_ptr[1:0] & 6'h4 == _io_out_weight_7_T_3[5:0] ? buffer_0_4 : _GEN_2310; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2312 = 2'h0 == read_ptr[1:0] & 6'h5 == _io_out_weight_7_T_3[5:0] ? buffer_0_5 : _GEN_2311; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2313 = 2'h0 == read_ptr[1:0] & 6'h6 == _io_out_weight_7_T_3[5:0] ? buffer_0_6 : _GEN_2312; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2314 = 2'h0 == read_ptr[1:0] & 6'h7 == _io_out_weight_7_T_3[5:0] ? buffer_0_7 : _GEN_2313; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2315 = 2'h0 == read_ptr[1:0] & 6'h8 == _io_out_weight_7_T_3[5:0] ? buffer_0_8 : _GEN_2314; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2316 = 2'h0 == read_ptr[1:0] & 6'h9 == _io_out_weight_7_T_3[5:0] ? buffer_0_9 : _GEN_2315; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2317 = 2'h0 == read_ptr[1:0] & 6'ha == _io_out_weight_7_T_3[5:0] ? buffer_0_10 : _GEN_2316; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2318 = 2'h0 == read_ptr[1:0] & 6'hb == _io_out_weight_7_T_3[5:0] ? buffer_0_11 : _GEN_2317; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2319 = 2'h0 == read_ptr[1:0] & 6'hc == _io_out_weight_7_T_3[5:0] ? buffer_0_12 : _GEN_2318; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2320 = 2'h0 == read_ptr[1:0] & 6'hd == _io_out_weight_7_T_3[5:0] ? buffer_0_13 : _GEN_2319; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2321 = 2'h0 == read_ptr[1:0] & 6'he == _io_out_weight_7_T_3[5:0] ? buffer_0_14 : _GEN_2320; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2322 = 2'h0 == read_ptr[1:0] & 6'hf == _io_out_weight_7_T_3[5:0] ? buffer_0_15 : _GEN_2321; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2323 = 2'h0 == read_ptr[1:0] & 6'h10 == _io_out_weight_7_T_3[5:0] ? buffer_0_16 : _GEN_2322; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2324 = 2'h0 == read_ptr[1:0] & 6'h11 == _io_out_weight_7_T_3[5:0] ? buffer_0_17 : _GEN_2323; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2325 = 2'h0 == read_ptr[1:0] & 6'h12 == _io_out_weight_7_T_3[5:0] ? buffer_0_18 : _GEN_2324; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2326 = 2'h0 == read_ptr[1:0] & 6'h13 == _io_out_weight_7_T_3[5:0] ? buffer_0_19 : _GEN_2325; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2327 = 2'h0 == read_ptr[1:0] & 6'h14 == _io_out_weight_7_T_3[5:0] ? buffer_0_20 : _GEN_2326; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2328 = 2'h0 == read_ptr[1:0] & 6'h15 == _io_out_weight_7_T_3[5:0] ? buffer_0_21 : _GEN_2327; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2329 = 2'h0 == read_ptr[1:0] & 6'h16 == _io_out_weight_7_T_3[5:0] ? buffer_0_22 : _GEN_2328; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2330 = 2'h0 == read_ptr[1:0] & 6'h17 == _io_out_weight_7_T_3[5:0] ? buffer_0_23 : _GEN_2329; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2331 = 2'h0 == read_ptr[1:0] & 6'h18 == _io_out_weight_7_T_3[5:0] ? buffer_0_24 : _GEN_2330; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2332 = 2'h0 == read_ptr[1:0] & 6'h19 == _io_out_weight_7_T_3[5:0] ? buffer_0_25 : _GEN_2331; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2333 = 2'h0 == read_ptr[1:0] & 6'h1a == _io_out_weight_7_T_3[5:0] ? buffer_0_26 : _GEN_2332; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2334 = 2'h0 == read_ptr[1:0] & 6'h1b == _io_out_weight_7_T_3[5:0] ? buffer_0_27 : _GEN_2333; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2335 = 2'h0 == read_ptr[1:0] & 6'h1c == _io_out_weight_7_T_3[5:0] ? buffer_0_28 : _GEN_2334; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2336 = 2'h0 == read_ptr[1:0] & 6'h1d == _io_out_weight_7_T_3[5:0] ? buffer_0_29 : _GEN_2335; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2337 = 2'h0 == read_ptr[1:0] & 6'h1e == _io_out_weight_7_T_3[5:0] ? buffer_0_30 : _GEN_2336; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2338 = 2'h0 == read_ptr[1:0] & 6'h1f == _io_out_weight_7_T_3[5:0] ? buffer_0_31 : _GEN_2337; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2339 = 2'h0 == read_ptr[1:0] & 6'h20 == _io_out_weight_7_T_3[5:0] ? buffer_0_32 : _GEN_2338; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2340 = 2'h0 == read_ptr[1:0] & 6'h21 == _io_out_weight_7_T_3[5:0] ? buffer_0_33 : _GEN_2339; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2341 = 2'h0 == read_ptr[1:0] & 6'h22 == _io_out_weight_7_T_3[5:0] ? buffer_0_34 : _GEN_2340; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2342 = 2'h0 == read_ptr[1:0] & 6'h23 == _io_out_weight_7_T_3[5:0] ? buffer_0_35 : _GEN_2341; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2343 = 2'h0 == read_ptr[1:0] & 6'h24 == _io_out_weight_7_T_3[5:0] ? buffer_0_36 : _GEN_2342; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2344 = 2'h0 == read_ptr[1:0] & 6'h25 == _io_out_weight_7_T_3[5:0] ? buffer_0_37 : _GEN_2343; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2345 = 2'h0 == read_ptr[1:0] & 6'h26 == _io_out_weight_7_T_3[5:0] ? buffer_0_38 : _GEN_2344; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2346 = 2'h0 == read_ptr[1:0] & 6'h27 == _io_out_weight_7_T_3[5:0] ? buffer_0_39 : _GEN_2345; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2347 = 2'h0 == read_ptr[1:0] & 6'h28 == _io_out_weight_7_T_3[5:0] ? buffer_0_40 : _GEN_2346; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2348 = 2'h0 == read_ptr[1:0] & 6'h29 == _io_out_weight_7_T_3[5:0] ? buffer_0_41 : _GEN_2347; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2349 = 2'h0 == read_ptr[1:0] & 6'h2a == _io_out_weight_7_T_3[5:0] ? buffer_0_42 : _GEN_2348; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2350 = 2'h0 == read_ptr[1:0] & 6'h2b == _io_out_weight_7_T_3[5:0] ? buffer_0_43 : _GEN_2349; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2351 = 2'h0 == read_ptr[1:0] & 6'h2c == _io_out_weight_7_T_3[5:0] ? buffer_0_44 : _GEN_2350; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2352 = 2'h0 == read_ptr[1:0] & 6'h2d == _io_out_weight_7_T_3[5:0] ? buffer_0_45 : _GEN_2351; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2353 = 2'h0 == read_ptr[1:0] & 6'h2e == _io_out_weight_7_T_3[5:0] ? buffer_0_46 : _GEN_2352; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2354 = 2'h0 == read_ptr[1:0] & 6'h2f == _io_out_weight_7_T_3[5:0] ? buffer_0_47 : _GEN_2353; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2355 = 2'h0 == read_ptr[1:0] & 6'h30 == _io_out_weight_7_T_3[5:0] ? buffer_0_48 : _GEN_2354; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2356 = 2'h0 == read_ptr[1:0] & 6'h31 == _io_out_weight_7_T_3[5:0] ? buffer_0_49 : _GEN_2355; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2357 = 2'h0 == read_ptr[1:0] & 6'h32 == _io_out_weight_7_T_3[5:0] ? buffer_0_50 : _GEN_2356; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2358 = 2'h0 == read_ptr[1:0] & 6'h33 == _io_out_weight_7_T_3[5:0] ? buffer_0_51 : _GEN_2357; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2359 = 2'h0 == read_ptr[1:0] & 6'h34 == _io_out_weight_7_T_3[5:0] ? buffer_0_52 : _GEN_2358; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2360 = 2'h0 == read_ptr[1:0] & 6'h35 == _io_out_weight_7_T_3[5:0] ? buffer_0_53 : _GEN_2359; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2361 = 2'h0 == read_ptr[1:0] & 6'h36 == _io_out_weight_7_T_3[5:0] ? buffer_0_54 : _GEN_2360; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2362 = 2'h0 == read_ptr[1:0] & 6'h37 == _io_out_weight_7_T_3[5:0] ? buffer_0_55 : _GEN_2361; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2363 = 2'h0 == read_ptr[1:0] & 6'h38 == _io_out_weight_7_T_3[5:0] ? buffer_0_56 : _GEN_2362; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2364 = 2'h0 == read_ptr[1:0] & 6'h39 == _io_out_weight_7_T_3[5:0] ? buffer_0_57 : _GEN_2363; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2365 = 2'h0 == read_ptr[1:0] & 6'h3a == _io_out_weight_7_T_3[5:0] ? buffer_0_58 : _GEN_2364; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2366 = 2'h0 == read_ptr[1:0] & 6'h3b == _io_out_weight_7_T_3[5:0] ? buffer_0_59 : _GEN_2365; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2367 = 2'h0 == read_ptr[1:0] & 6'h3c == _io_out_weight_7_T_3[5:0] ? buffer_0_60 : _GEN_2366; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2368 = 2'h0 == read_ptr[1:0] & 6'h3d == _io_out_weight_7_T_3[5:0] ? buffer_0_61 : _GEN_2367; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2369 = 2'h0 == read_ptr[1:0] & 6'h3e == _io_out_weight_7_T_3[5:0] ? buffer_0_62 : _GEN_2368; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2370 = 2'h0 == read_ptr[1:0] & 6'h3f == _io_out_weight_7_T_3[5:0] ? buffer_0_63 : _GEN_2369; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2371 = 2'h1 == read_ptr[1:0] & 6'h0 == _io_out_weight_7_T_3[5:0] ? buffer_1_0 : _GEN_2370; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2372 = 2'h1 == read_ptr[1:0] & 6'h1 == _io_out_weight_7_T_3[5:0] ? buffer_1_1 : _GEN_2371; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2373 = 2'h1 == read_ptr[1:0] & 6'h2 == _io_out_weight_7_T_3[5:0] ? buffer_1_2 : _GEN_2372; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2374 = 2'h1 == read_ptr[1:0] & 6'h3 == _io_out_weight_7_T_3[5:0] ? buffer_1_3 : _GEN_2373; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2375 = 2'h1 == read_ptr[1:0] & 6'h4 == _io_out_weight_7_T_3[5:0] ? buffer_1_4 : _GEN_2374; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2376 = 2'h1 == read_ptr[1:0] & 6'h5 == _io_out_weight_7_T_3[5:0] ? buffer_1_5 : _GEN_2375; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2377 = 2'h1 == read_ptr[1:0] & 6'h6 == _io_out_weight_7_T_3[5:0] ? buffer_1_6 : _GEN_2376; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2378 = 2'h1 == read_ptr[1:0] & 6'h7 == _io_out_weight_7_T_3[5:0] ? buffer_1_7 : _GEN_2377; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2379 = 2'h1 == read_ptr[1:0] & 6'h8 == _io_out_weight_7_T_3[5:0] ? buffer_1_8 : _GEN_2378; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2380 = 2'h1 == read_ptr[1:0] & 6'h9 == _io_out_weight_7_T_3[5:0] ? buffer_1_9 : _GEN_2379; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2381 = 2'h1 == read_ptr[1:0] & 6'ha == _io_out_weight_7_T_3[5:0] ? buffer_1_10 : _GEN_2380; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2382 = 2'h1 == read_ptr[1:0] & 6'hb == _io_out_weight_7_T_3[5:0] ? buffer_1_11 : _GEN_2381; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2383 = 2'h1 == read_ptr[1:0] & 6'hc == _io_out_weight_7_T_3[5:0] ? buffer_1_12 : _GEN_2382; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2384 = 2'h1 == read_ptr[1:0] & 6'hd == _io_out_weight_7_T_3[5:0] ? buffer_1_13 : _GEN_2383; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2385 = 2'h1 == read_ptr[1:0] & 6'he == _io_out_weight_7_T_3[5:0] ? buffer_1_14 : _GEN_2384; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2386 = 2'h1 == read_ptr[1:0] & 6'hf == _io_out_weight_7_T_3[5:0] ? buffer_1_15 : _GEN_2385; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2387 = 2'h1 == read_ptr[1:0] & 6'h10 == _io_out_weight_7_T_3[5:0] ? buffer_1_16 : _GEN_2386; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2388 = 2'h1 == read_ptr[1:0] & 6'h11 == _io_out_weight_7_T_3[5:0] ? buffer_1_17 : _GEN_2387; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2389 = 2'h1 == read_ptr[1:0] & 6'h12 == _io_out_weight_7_T_3[5:0] ? buffer_1_18 : _GEN_2388; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2390 = 2'h1 == read_ptr[1:0] & 6'h13 == _io_out_weight_7_T_3[5:0] ? buffer_1_19 : _GEN_2389; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2391 = 2'h1 == read_ptr[1:0] & 6'h14 == _io_out_weight_7_T_3[5:0] ? buffer_1_20 : _GEN_2390; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2392 = 2'h1 == read_ptr[1:0] & 6'h15 == _io_out_weight_7_T_3[5:0] ? buffer_1_21 : _GEN_2391; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2393 = 2'h1 == read_ptr[1:0] & 6'h16 == _io_out_weight_7_T_3[5:0] ? buffer_1_22 : _GEN_2392; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2394 = 2'h1 == read_ptr[1:0] & 6'h17 == _io_out_weight_7_T_3[5:0] ? buffer_1_23 : _GEN_2393; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2395 = 2'h1 == read_ptr[1:0] & 6'h18 == _io_out_weight_7_T_3[5:0] ? buffer_1_24 : _GEN_2394; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2396 = 2'h1 == read_ptr[1:0] & 6'h19 == _io_out_weight_7_T_3[5:0] ? buffer_1_25 : _GEN_2395; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2397 = 2'h1 == read_ptr[1:0] & 6'h1a == _io_out_weight_7_T_3[5:0] ? buffer_1_26 : _GEN_2396; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2398 = 2'h1 == read_ptr[1:0] & 6'h1b == _io_out_weight_7_T_3[5:0] ? buffer_1_27 : _GEN_2397; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2399 = 2'h1 == read_ptr[1:0] & 6'h1c == _io_out_weight_7_T_3[5:0] ? buffer_1_28 : _GEN_2398; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2400 = 2'h1 == read_ptr[1:0] & 6'h1d == _io_out_weight_7_T_3[5:0] ? buffer_1_29 : _GEN_2399; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2401 = 2'h1 == read_ptr[1:0] & 6'h1e == _io_out_weight_7_T_3[5:0] ? buffer_1_30 : _GEN_2400; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2402 = 2'h1 == read_ptr[1:0] & 6'h1f == _io_out_weight_7_T_3[5:0] ? buffer_1_31 : _GEN_2401; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2403 = 2'h1 == read_ptr[1:0] & 6'h20 == _io_out_weight_7_T_3[5:0] ? buffer_1_32 : _GEN_2402; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2404 = 2'h1 == read_ptr[1:0] & 6'h21 == _io_out_weight_7_T_3[5:0] ? buffer_1_33 : _GEN_2403; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2405 = 2'h1 == read_ptr[1:0] & 6'h22 == _io_out_weight_7_T_3[5:0] ? buffer_1_34 : _GEN_2404; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2406 = 2'h1 == read_ptr[1:0] & 6'h23 == _io_out_weight_7_T_3[5:0] ? buffer_1_35 : _GEN_2405; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2407 = 2'h1 == read_ptr[1:0] & 6'h24 == _io_out_weight_7_T_3[5:0] ? buffer_1_36 : _GEN_2406; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2408 = 2'h1 == read_ptr[1:0] & 6'h25 == _io_out_weight_7_T_3[5:0] ? buffer_1_37 : _GEN_2407; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2409 = 2'h1 == read_ptr[1:0] & 6'h26 == _io_out_weight_7_T_3[5:0] ? buffer_1_38 : _GEN_2408; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2410 = 2'h1 == read_ptr[1:0] & 6'h27 == _io_out_weight_7_T_3[5:0] ? buffer_1_39 : _GEN_2409; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2411 = 2'h1 == read_ptr[1:0] & 6'h28 == _io_out_weight_7_T_3[5:0] ? buffer_1_40 : _GEN_2410; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2412 = 2'h1 == read_ptr[1:0] & 6'h29 == _io_out_weight_7_T_3[5:0] ? buffer_1_41 : _GEN_2411; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2413 = 2'h1 == read_ptr[1:0] & 6'h2a == _io_out_weight_7_T_3[5:0] ? buffer_1_42 : _GEN_2412; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2414 = 2'h1 == read_ptr[1:0] & 6'h2b == _io_out_weight_7_T_3[5:0] ? buffer_1_43 : _GEN_2413; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2415 = 2'h1 == read_ptr[1:0] & 6'h2c == _io_out_weight_7_T_3[5:0] ? buffer_1_44 : _GEN_2414; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2416 = 2'h1 == read_ptr[1:0] & 6'h2d == _io_out_weight_7_T_3[5:0] ? buffer_1_45 : _GEN_2415; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2417 = 2'h1 == read_ptr[1:0] & 6'h2e == _io_out_weight_7_T_3[5:0] ? buffer_1_46 : _GEN_2416; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2418 = 2'h1 == read_ptr[1:0] & 6'h2f == _io_out_weight_7_T_3[5:0] ? buffer_1_47 : _GEN_2417; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2419 = 2'h1 == read_ptr[1:0] & 6'h30 == _io_out_weight_7_T_3[5:0] ? buffer_1_48 : _GEN_2418; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2420 = 2'h1 == read_ptr[1:0] & 6'h31 == _io_out_weight_7_T_3[5:0] ? buffer_1_49 : _GEN_2419; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2421 = 2'h1 == read_ptr[1:0] & 6'h32 == _io_out_weight_7_T_3[5:0] ? buffer_1_50 : _GEN_2420; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2422 = 2'h1 == read_ptr[1:0] & 6'h33 == _io_out_weight_7_T_3[5:0] ? buffer_1_51 : _GEN_2421; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2423 = 2'h1 == read_ptr[1:0] & 6'h34 == _io_out_weight_7_T_3[5:0] ? buffer_1_52 : _GEN_2422; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2424 = 2'h1 == read_ptr[1:0] & 6'h35 == _io_out_weight_7_T_3[5:0] ? buffer_1_53 : _GEN_2423; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2425 = 2'h1 == read_ptr[1:0] & 6'h36 == _io_out_weight_7_T_3[5:0] ? buffer_1_54 : _GEN_2424; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2426 = 2'h1 == read_ptr[1:0] & 6'h37 == _io_out_weight_7_T_3[5:0] ? buffer_1_55 : _GEN_2425; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2427 = 2'h1 == read_ptr[1:0] & 6'h38 == _io_out_weight_7_T_3[5:0] ? buffer_1_56 : _GEN_2426; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2428 = 2'h1 == read_ptr[1:0] & 6'h39 == _io_out_weight_7_T_3[5:0] ? buffer_1_57 : _GEN_2427; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2429 = 2'h1 == read_ptr[1:0] & 6'h3a == _io_out_weight_7_T_3[5:0] ? buffer_1_58 : _GEN_2428; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2430 = 2'h1 == read_ptr[1:0] & 6'h3b == _io_out_weight_7_T_3[5:0] ? buffer_1_59 : _GEN_2429; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2431 = 2'h1 == read_ptr[1:0] & 6'h3c == _io_out_weight_7_T_3[5:0] ? buffer_1_60 : _GEN_2430; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2432 = 2'h1 == read_ptr[1:0] & 6'h3d == _io_out_weight_7_T_3[5:0] ? buffer_1_61 : _GEN_2431; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2433 = 2'h1 == read_ptr[1:0] & 6'h3e == _io_out_weight_7_T_3[5:0] ? buffer_1_62 : _GEN_2432; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2434 = 2'h1 == read_ptr[1:0] & 6'h3f == _io_out_weight_7_T_3[5:0] ? buffer_1_63 : _GEN_2433; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2435 = 2'h2 == read_ptr[1:0] & 6'h0 == _io_out_weight_7_T_3[5:0] ? buffer_2_0 : _GEN_2434; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2436 = 2'h2 == read_ptr[1:0] & 6'h1 == _io_out_weight_7_T_3[5:0] ? buffer_2_1 : _GEN_2435; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2437 = 2'h2 == read_ptr[1:0] & 6'h2 == _io_out_weight_7_T_3[5:0] ? buffer_2_2 : _GEN_2436; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2438 = 2'h2 == read_ptr[1:0] & 6'h3 == _io_out_weight_7_T_3[5:0] ? buffer_2_3 : _GEN_2437; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2439 = 2'h2 == read_ptr[1:0] & 6'h4 == _io_out_weight_7_T_3[5:0] ? buffer_2_4 : _GEN_2438; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2440 = 2'h2 == read_ptr[1:0] & 6'h5 == _io_out_weight_7_T_3[5:0] ? buffer_2_5 : _GEN_2439; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2441 = 2'h2 == read_ptr[1:0] & 6'h6 == _io_out_weight_7_T_3[5:0] ? buffer_2_6 : _GEN_2440; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2442 = 2'h2 == read_ptr[1:0] & 6'h7 == _io_out_weight_7_T_3[5:0] ? buffer_2_7 : _GEN_2441; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2443 = 2'h2 == read_ptr[1:0] & 6'h8 == _io_out_weight_7_T_3[5:0] ? buffer_2_8 : _GEN_2442; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2444 = 2'h2 == read_ptr[1:0] & 6'h9 == _io_out_weight_7_T_3[5:0] ? buffer_2_9 : _GEN_2443; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2445 = 2'h2 == read_ptr[1:0] & 6'ha == _io_out_weight_7_T_3[5:0] ? buffer_2_10 : _GEN_2444; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2446 = 2'h2 == read_ptr[1:0] & 6'hb == _io_out_weight_7_T_3[5:0] ? buffer_2_11 : _GEN_2445; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2447 = 2'h2 == read_ptr[1:0] & 6'hc == _io_out_weight_7_T_3[5:0] ? buffer_2_12 : _GEN_2446; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2448 = 2'h2 == read_ptr[1:0] & 6'hd == _io_out_weight_7_T_3[5:0] ? buffer_2_13 : _GEN_2447; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2449 = 2'h2 == read_ptr[1:0] & 6'he == _io_out_weight_7_T_3[5:0] ? buffer_2_14 : _GEN_2448; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2450 = 2'h2 == read_ptr[1:0] & 6'hf == _io_out_weight_7_T_3[5:0] ? buffer_2_15 : _GEN_2449; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2451 = 2'h2 == read_ptr[1:0] & 6'h10 == _io_out_weight_7_T_3[5:0] ? buffer_2_16 : _GEN_2450; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2452 = 2'h2 == read_ptr[1:0] & 6'h11 == _io_out_weight_7_T_3[5:0] ? buffer_2_17 : _GEN_2451; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2453 = 2'h2 == read_ptr[1:0] & 6'h12 == _io_out_weight_7_T_3[5:0] ? buffer_2_18 : _GEN_2452; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2454 = 2'h2 == read_ptr[1:0] & 6'h13 == _io_out_weight_7_T_3[5:0] ? buffer_2_19 : _GEN_2453; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2455 = 2'h2 == read_ptr[1:0] & 6'h14 == _io_out_weight_7_T_3[5:0] ? buffer_2_20 : _GEN_2454; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2456 = 2'h2 == read_ptr[1:0] & 6'h15 == _io_out_weight_7_T_3[5:0] ? buffer_2_21 : _GEN_2455; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2457 = 2'h2 == read_ptr[1:0] & 6'h16 == _io_out_weight_7_T_3[5:0] ? buffer_2_22 : _GEN_2456; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2458 = 2'h2 == read_ptr[1:0] & 6'h17 == _io_out_weight_7_T_3[5:0] ? buffer_2_23 : _GEN_2457; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2459 = 2'h2 == read_ptr[1:0] & 6'h18 == _io_out_weight_7_T_3[5:0] ? buffer_2_24 : _GEN_2458; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2460 = 2'h2 == read_ptr[1:0] & 6'h19 == _io_out_weight_7_T_3[5:0] ? buffer_2_25 : _GEN_2459; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2461 = 2'h2 == read_ptr[1:0] & 6'h1a == _io_out_weight_7_T_3[5:0] ? buffer_2_26 : _GEN_2460; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2462 = 2'h2 == read_ptr[1:0] & 6'h1b == _io_out_weight_7_T_3[5:0] ? buffer_2_27 : _GEN_2461; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2463 = 2'h2 == read_ptr[1:0] & 6'h1c == _io_out_weight_7_T_3[5:0] ? buffer_2_28 : _GEN_2462; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2464 = 2'h2 == read_ptr[1:0] & 6'h1d == _io_out_weight_7_T_3[5:0] ? buffer_2_29 : _GEN_2463; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2465 = 2'h2 == read_ptr[1:0] & 6'h1e == _io_out_weight_7_T_3[5:0] ? buffer_2_30 : _GEN_2464; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2466 = 2'h2 == read_ptr[1:0] & 6'h1f == _io_out_weight_7_T_3[5:0] ? buffer_2_31 : _GEN_2465; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2467 = 2'h2 == read_ptr[1:0] & 6'h20 == _io_out_weight_7_T_3[5:0] ? buffer_2_32 : _GEN_2466; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2468 = 2'h2 == read_ptr[1:0] & 6'h21 == _io_out_weight_7_T_3[5:0] ? buffer_2_33 : _GEN_2467; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2469 = 2'h2 == read_ptr[1:0] & 6'h22 == _io_out_weight_7_T_3[5:0] ? buffer_2_34 : _GEN_2468; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2470 = 2'h2 == read_ptr[1:0] & 6'h23 == _io_out_weight_7_T_3[5:0] ? buffer_2_35 : _GEN_2469; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2471 = 2'h2 == read_ptr[1:0] & 6'h24 == _io_out_weight_7_T_3[5:0] ? buffer_2_36 : _GEN_2470; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2472 = 2'h2 == read_ptr[1:0] & 6'h25 == _io_out_weight_7_T_3[5:0] ? buffer_2_37 : _GEN_2471; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2473 = 2'h2 == read_ptr[1:0] & 6'h26 == _io_out_weight_7_T_3[5:0] ? buffer_2_38 : _GEN_2472; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2474 = 2'h2 == read_ptr[1:0] & 6'h27 == _io_out_weight_7_T_3[5:0] ? buffer_2_39 : _GEN_2473; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2475 = 2'h2 == read_ptr[1:0] & 6'h28 == _io_out_weight_7_T_3[5:0] ? buffer_2_40 : _GEN_2474; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2476 = 2'h2 == read_ptr[1:0] & 6'h29 == _io_out_weight_7_T_3[5:0] ? buffer_2_41 : _GEN_2475; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2477 = 2'h2 == read_ptr[1:0] & 6'h2a == _io_out_weight_7_T_3[5:0] ? buffer_2_42 : _GEN_2476; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2478 = 2'h2 == read_ptr[1:0] & 6'h2b == _io_out_weight_7_T_3[5:0] ? buffer_2_43 : _GEN_2477; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2479 = 2'h2 == read_ptr[1:0] & 6'h2c == _io_out_weight_7_T_3[5:0] ? buffer_2_44 : _GEN_2478; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2480 = 2'h2 == read_ptr[1:0] & 6'h2d == _io_out_weight_7_T_3[5:0] ? buffer_2_45 : _GEN_2479; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2481 = 2'h2 == read_ptr[1:0] & 6'h2e == _io_out_weight_7_T_3[5:0] ? buffer_2_46 : _GEN_2480; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2482 = 2'h2 == read_ptr[1:0] & 6'h2f == _io_out_weight_7_T_3[5:0] ? buffer_2_47 : _GEN_2481; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2483 = 2'h2 == read_ptr[1:0] & 6'h30 == _io_out_weight_7_T_3[5:0] ? buffer_2_48 : _GEN_2482; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2484 = 2'h2 == read_ptr[1:0] & 6'h31 == _io_out_weight_7_T_3[5:0] ? buffer_2_49 : _GEN_2483; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2485 = 2'h2 == read_ptr[1:0] & 6'h32 == _io_out_weight_7_T_3[5:0] ? buffer_2_50 : _GEN_2484; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2486 = 2'h2 == read_ptr[1:0] & 6'h33 == _io_out_weight_7_T_3[5:0] ? buffer_2_51 : _GEN_2485; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2487 = 2'h2 == read_ptr[1:0] & 6'h34 == _io_out_weight_7_T_3[5:0] ? buffer_2_52 : _GEN_2486; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2488 = 2'h2 == read_ptr[1:0] & 6'h35 == _io_out_weight_7_T_3[5:0] ? buffer_2_53 : _GEN_2487; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2489 = 2'h2 == read_ptr[1:0] & 6'h36 == _io_out_weight_7_T_3[5:0] ? buffer_2_54 : _GEN_2488; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2490 = 2'h2 == read_ptr[1:0] & 6'h37 == _io_out_weight_7_T_3[5:0] ? buffer_2_55 : _GEN_2489; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2491 = 2'h2 == read_ptr[1:0] & 6'h38 == _io_out_weight_7_T_3[5:0] ? buffer_2_56 : _GEN_2490; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2492 = 2'h2 == read_ptr[1:0] & 6'h39 == _io_out_weight_7_T_3[5:0] ? buffer_2_57 : _GEN_2491; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2493 = 2'h2 == read_ptr[1:0] & 6'h3a == _io_out_weight_7_T_3[5:0] ? buffer_2_58 : _GEN_2492; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2494 = 2'h2 == read_ptr[1:0] & 6'h3b == _io_out_weight_7_T_3[5:0] ? buffer_2_59 : _GEN_2493; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2495 = 2'h2 == read_ptr[1:0] & 6'h3c == _io_out_weight_7_T_3[5:0] ? buffer_2_60 : _GEN_2494; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2496 = 2'h2 == read_ptr[1:0] & 6'h3d == _io_out_weight_7_T_3[5:0] ? buffer_2_61 : _GEN_2495; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2497 = 2'h2 == read_ptr[1:0] & 6'h3e == _io_out_weight_7_T_3[5:0] ? buffer_2_62 : _GEN_2496; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2498 = 2'h2 == read_ptr[1:0] & 6'h3f == _io_out_weight_7_T_3[5:0] ? buffer_2_63 : _GEN_2497; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2499 = 2'h3 == read_ptr[1:0] & 6'h0 == _io_out_weight_7_T_3[5:0] ? buffer_3_0 : _GEN_2498; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2500 = 2'h3 == read_ptr[1:0] & 6'h1 == _io_out_weight_7_T_3[5:0] ? buffer_3_1 : _GEN_2499; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2501 = 2'h3 == read_ptr[1:0] & 6'h2 == _io_out_weight_7_T_3[5:0] ? buffer_3_2 : _GEN_2500; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2502 = 2'h3 == read_ptr[1:0] & 6'h3 == _io_out_weight_7_T_3[5:0] ? buffer_3_3 : _GEN_2501; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2503 = 2'h3 == read_ptr[1:0] & 6'h4 == _io_out_weight_7_T_3[5:0] ? buffer_3_4 : _GEN_2502; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2504 = 2'h3 == read_ptr[1:0] & 6'h5 == _io_out_weight_7_T_3[5:0] ? buffer_3_5 : _GEN_2503; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2505 = 2'h3 == read_ptr[1:0] & 6'h6 == _io_out_weight_7_T_3[5:0] ? buffer_3_6 : _GEN_2504; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2506 = 2'h3 == read_ptr[1:0] & 6'h7 == _io_out_weight_7_T_3[5:0] ? buffer_3_7 : _GEN_2505; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2507 = 2'h3 == read_ptr[1:0] & 6'h8 == _io_out_weight_7_T_3[5:0] ? buffer_3_8 : _GEN_2506; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2508 = 2'h3 == read_ptr[1:0] & 6'h9 == _io_out_weight_7_T_3[5:0] ? buffer_3_9 : _GEN_2507; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2509 = 2'h3 == read_ptr[1:0] & 6'ha == _io_out_weight_7_T_3[5:0] ? buffer_3_10 : _GEN_2508; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2510 = 2'h3 == read_ptr[1:0] & 6'hb == _io_out_weight_7_T_3[5:0] ? buffer_3_11 : _GEN_2509; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2511 = 2'h3 == read_ptr[1:0] & 6'hc == _io_out_weight_7_T_3[5:0] ? buffer_3_12 : _GEN_2510; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2512 = 2'h3 == read_ptr[1:0] & 6'hd == _io_out_weight_7_T_3[5:0] ? buffer_3_13 : _GEN_2511; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2513 = 2'h3 == read_ptr[1:0] & 6'he == _io_out_weight_7_T_3[5:0] ? buffer_3_14 : _GEN_2512; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2514 = 2'h3 == read_ptr[1:0] & 6'hf == _io_out_weight_7_T_3[5:0] ? buffer_3_15 : _GEN_2513; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2515 = 2'h3 == read_ptr[1:0] & 6'h10 == _io_out_weight_7_T_3[5:0] ? buffer_3_16 : _GEN_2514; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2516 = 2'h3 == read_ptr[1:0] & 6'h11 == _io_out_weight_7_T_3[5:0] ? buffer_3_17 : _GEN_2515; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2517 = 2'h3 == read_ptr[1:0] & 6'h12 == _io_out_weight_7_T_3[5:0] ? buffer_3_18 : _GEN_2516; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2518 = 2'h3 == read_ptr[1:0] & 6'h13 == _io_out_weight_7_T_3[5:0] ? buffer_3_19 : _GEN_2517; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2519 = 2'h3 == read_ptr[1:0] & 6'h14 == _io_out_weight_7_T_3[5:0] ? buffer_3_20 : _GEN_2518; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2520 = 2'h3 == read_ptr[1:0] & 6'h15 == _io_out_weight_7_T_3[5:0] ? buffer_3_21 : _GEN_2519; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2521 = 2'h3 == read_ptr[1:0] & 6'h16 == _io_out_weight_7_T_3[5:0] ? buffer_3_22 : _GEN_2520; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2522 = 2'h3 == read_ptr[1:0] & 6'h17 == _io_out_weight_7_T_3[5:0] ? buffer_3_23 : _GEN_2521; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2523 = 2'h3 == read_ptr[1:0] & 6'h18 == _io_out_weight_7_T_3[5:0] ? buffer_3_24 : _GEN_2522; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2524 = 2'h3 == read_ptr[1:0] & 6'h19 == _io_out_weight_7_T_3[5:0] ? buffer_3_25 : _GEN_2523; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2525 = 2'h3 == read_ptr[1:0] & 6'h1a == _io_out_weight_7_T_3[5:0] ? buffer_3_26 : _GEN_2524; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2526 = 2'h3 == read_ptr[1:0] & 6'h1b == _io_out_weight_7_T_3[5:0] ? buffer_3_27 : _GEN_2525; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2527 = 2'h3 == read_ptr[1:0] & 6'h1c == _io_out_weight_7_T_3[5:0] ? buffer_3_28 : _GEN_2526; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2528 = 2'h3 == read_ptr[1:0] & 6'h1d == _io_out_weight_7_T_3[5:0] ? buffer_3_29 : _GEN_2527; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2529 = 2'h3 == read_ptr[1:0] & 6'h1e == _io_out_weight_7_T_3[5:0] ? buffer_3_30 : _GEN_2528; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2530 = 2'h3 == read_ptr[1:0] & 6'h1f == _io_out_weight_7_T_3[5:0] ? buffer_3_31 : _GEN_2529; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2531 = 2'h3 == read_ptr[1:0] & 6'h20 == _io_out_weight_7_T_3[5:0] ? buffer_3_32 : _GEN_2530; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2532 = 2'h3 == read_ptr[1:0] & 6'h21 == _io_out_weight_7_T_3[5:0] ? buffer_3_33 : _GEN_2531; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2533 = 2'h3 == read_ptr[1:0] & 6'h22 == _io_out_weight_7_T_3[5:0] ? buffer_3_34 : _GEN_2532; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2534 = 2'h3 == read_ptr[1:0] & 6'h23 == _io_out_weight_7_T_3[5:0] ? buffer_3_35 : _GEN_2533; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2535 = 2'h3 == read_ptr[1:0] & 6'h24 == _io_out_weight_7_T_3[5:0] ? buffer_3_36 : _GEN_2534; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2536 = 2'h3 == read_ptr[1:0] & 6'h25 == _io_out_weight_7_T_3[5:0] ? buffer_3_37 : _GEN_2535; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2537 = 2'h3 == read_ptr[1:0] & 6'h26 == _io_out_weight_7_T_3[5:0] ? buffer_3_38 : _GEN_2536; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2538 = 2'h3 == read_ptr[1:0] & 6'h27 == _io_out_weight_7_T_3[5:0] ? buffer_3_39 : _GEN_2537; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2539 = 2'h3 == read_ptr[1:0] & 6'h28 == _io_out_weight_7_T_3[5:0] ? buffer_3_40 : _GEN_2538; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2540 = 2'h3 == read_ptr[1:0] & 6'h29 == _io_out_weight_7_T_3[5:0] ? buffer_3_41 : _GEN_2539; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2541 = 2'h3 == read_ptr[1:0] & 6'h2a == _io_out_weight_7_T_3[5:0] ? buffer_3_42 : _GEN_2540; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2542 = 2'h3 == read_ptr[1:0] & 6'h2b == _io_out_weight_7_T_3[5:0] ? buffer_3_43 : _GEN_2541; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2543 = 2'h3 == read_ptr[1:0] & 6'h2c == _io_out_weight_7_T_3[5:0] ? buffer_3_44 : _GEN_2542; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2544 = 2'h3 == read_ptr[1:0] & 6'h2d == _io_out_weight_7_T_3[5:0] ? buffer_3_45 : _GEN_2543; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2545 = 2'h3 == read_ptr[1:0] & 6'h2e == _io_out_weight_7_T_3[5:0] ? buffer_3_46 : _GEN_2544; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2546 = 2'h3 == read_ptr[1:0] & 6'h2f == _io_out_weight_7_T_3[5:0] ? buffer_3_47 : _GEN_2545; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2547 = 2'h3 == read_ptr[1:0] & 6'h30 == _io_out_weight_7_T_3[5:0] ? buffer_3_48 : _GEN_2546; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2548 = 2'h3 == read_ptr[1:0] & 6'h31 == _io_out_weight_7_T_3[5:0] ? buffer_3_49 : _GEN_2547; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2549 = 2'h3 == read_ptr[1:0] & 6'h32 == _io_out_weight_7_T_3[5:0] ? buffer_3_50 : _GEN_2548; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2550 = 2'h3 == read_ptr[1:0] & 6'h33 == _io_out_weight_7_T_3[5:0] ? buffer_3_51 : _GEN_2549; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2551 = 2'h3 == read_ptr[1:0] & 6'h34 == _io_out_weight_7_T_3[5:0] ? buffer_3_52 : _GEN_2550; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2552 = 2'h3 == read_ptr[1:0] & 6'h35 == _io_out_weight_7_T_3[5:0] ? buffer_3_53 : _GEN_2551; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2553 = 2'h3 == read_ptr[1:0] & 6'h36 == _io_out_weight_7_T_3[5:0] ? buffer_3_54 : _GEN_2552; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2554 = 2'h3 == read_ptr[1:0] & 6'h37 == _io_out_weight_7_T_3[5:0] ? buffer_3_55 : _GEN_2553; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2555 = 2'h3 == read_ptr[1:0] & 6'h38 == _io_out_weight_7_T_3[5:0] ? buffer_3_56 : _GEN_2554; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2556 = 2'h3 == read_ptr[1:0] & 6'h39 == _io_out_weight_7_T_3[5:0] ? buffer_3_57 : _GEN_2555; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2557 = 2'h3 == read_ptr[1:0] & 6'h3a == _io_out_weight_7_T_3[5:0] ? buffer_3_58 : _GEN_2556; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2558 = 2'h3 == read_ptr[1:0] & 6'h3b == _io_out_weight_7_T_3[5:0] ? buffer_3_59 : _GEN_2557; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2559 = 2'h3 == read_ptr[1:0] & 6'h3c == _io_out_weight_7_T_3[5:0] ? buffer_3_60 : _GEN_2558; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2560 = 2'h3 == read_ptr[1:0] & 6'h3d == _io_out_weight_7_T_3[5:0] ? buffer_3_61 : _GEN_2559; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2561 = 2'h3 == read_ptr[1:0] & 6'h3e == _io_out_weight_7_T_3[5:0] ? buffer_3_62 : _GEN_2560; // @[Weight_Buffer.scala 64:{24,24}]
  wire [7:0] _GEN_2562 = 2'h3 == read_ptr[1:0] & 6'h3f == _io_out_weight_7_T_3[5:0] ? buffer_3_63 : _GEN_2561; // @[Weight_Buffer.scala 64:{24,24}]
  wire [2:0] _read_ptr_T_1 = read_ptr + 3'h1; // @[Weight_Buffer.scala 74:26]
  assign io_out_weight_0 = shift_ptr != 4'h8 ? _GEN_770 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_1 = shift_ptr != 4'h8 ? _GEN_1026 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_2 = shift_ptr != 4'h8 ? _GEN_1282 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_3 = shift_ptr != 4'h8 ? _GEN_1538 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_4 = shift_ptr != 4'h8 ? _GEN_1794 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_5 = shift_ptr != 4'h8 ? _GEN_2050 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_6 = shift_ptr != 4'h8 ? _GEN_2306 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_weight_7 = shift_ptr != 4'h8 ? _GEN_2562 : 8'h0; // @[Weight_Buffer.scala 61:34 64:24 69:24]
  assign io_out_shift = shift_ptr != 4'h8; // @[Weight_Buffer.scala 61:18]
  assign io_isfull = read_ptr[1:0] == write_ptr[1:0] & read_ptr[2] != write_ptr[2]; // @[Weight_Buffer.scala 34:78]
  assign io_isempty = _full_T_2 & read_ptr[2] == write_ptr[2]; // @[Weight_Buffer.scala 35:79]
  assign io_isdone = shift_ptr == 4'h0; // @[Weight_Buffer.scala 79:18]
  always @(posedge clock) begin
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_0 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_0 <= io_in_weight_x_0; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_1 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_1 <= io_in_weight_x_1; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_2 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_2 <= io_in_weight_x_2; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_3 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_3 <= io_in_weight_x_3; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_4 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_4 <= io_in_weight_x_4; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_5 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_5 <= io_in_weight_x_5; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_6 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_6 <= io_in_weight_x_6; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_7 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_7 <= io_in_weight_x_7; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_8 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_8 <= io_in_weight_x_8; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_9 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_9 <= io_in_weight_x_9; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_10 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_10 <= io_in_weight_x_10; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_11 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_11 <= io_in_weight_x_11; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_12 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_12 <= io_in_weight_x_12; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_13 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_13 <= io_in_weight_x_13; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_14 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_14 <= io_in_weight_x_14; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_15 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_15 <= io_in_weight_x_15; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_16 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_16 <= io_in_weight_x_16; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_17 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_17 <= io_in_weight_x_17; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_18 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_18 <= io_in_weight_x_18; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_19 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_19 <= io_in_weight_x_19; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_20 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_20 <= io_in_weight_x_20; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_21 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_21 <= io_in_weight_x_21; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_22 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_22 <= io_in_weight_x_22; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_23 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_23 <= io_in_weight_x_23; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_24 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_24 <= io_in_weight_x_24; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_25 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_25 <= io_in_weight_x_25; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_26 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_26 <= io_in_weight_x_26; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_27 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_27 <= io_in_weight_x_27; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_28 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_28 <= io_in_weight_x_28; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_29 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_29 <= io_in_weight_x_29; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_30 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_30 <= io_in_weight_x_30; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_31 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_31 <= io_in_weight_x_31; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_32 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_32 <= io_in_weight_x_32; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_33 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_33 <= io_in_weight_x_33; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_34 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_34 <= io_in_weight_x_34; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_35 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_35 <= io_in_weight_x_35; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_36 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_36 <= io_in_weight_x_36; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_37 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_37 <= io_in_weight_x_37; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_38 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_38 <= io_in_weight_x_38; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_39 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_39 <= io_in_weight_x_39; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_40 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_40 <= io_in_weight_x_40; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_41 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_41 <= io_in_weight_x_41; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_42 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_42 <= io_in_weight_x_42; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_43 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_43 <= io_in_weight_x_43; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_44 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_44 <= io_in_weight_x_44; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_45 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_45 <= io_in_weight_x_45; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_46 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_46 <= io_in_weight_x_46; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_47 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_47 <= io_in_weight_x_47; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_48 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_48 <= io_in_weight_x_48; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_49 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_49 <= io_in_weight_x_49; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_50 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_50 <= io_in_weight_x_50; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_51 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_51 <= io_in_weight_x_51; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_52 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_52 <= io_in_weight_x_52; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_53 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_53 <= io_in_weight_x_53; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_54 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_54 <= io_in_weight_x_54; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_55 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_55 <= io_in_weight_x_55; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_56 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_56 <= io_in_weight_x_56; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_57 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_57 <= io_in_weight_x_57; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_58 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_58 <= io_in_weight_x_58; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_59 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_59 <= io_in_weight_x_59; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_60 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_60 <= io_in_weight_x_60; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_61 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_61 <= io_in_weight_x_61; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_62 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_62 <= io_in_weight_x_62; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_0_63 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h0 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_0_63 <= io_in_weight_x_63; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_0 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_0 <= io_in_weight_x_0; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_1 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_1 <= io_in_weight_x_1; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_2 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_2 <= io_in_weight_x_2; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_3 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_3 <= io_in_weight_x_3; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_4 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_4 <= io_in_weight_x_4; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_5 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_5 <= io_in_weight_x_5; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_6 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_6 <= io_in_weight_x_6; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_7 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_7 <= io_in_weight_x_7; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_8 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_8 <= io_in_weight_x_8; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_9 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_9 <= io_in_weight_x_9; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_10 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_10 <= io_in_weight_x_10; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_11 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_11 <= io_in_weight_x_11; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_12 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_12 <= io_in_weight_x_12; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_13 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_13 <= io_in_weight_x_13; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_14 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_14 <= io_in_weight_x_14; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_15 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_15 <= io_in_weight_x_15; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_16 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_16 <= io_in_weight_x_16; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_17 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_17 <= io_in_weight_x_17; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_18 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_18 <= io_in_weight_x_18; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_19 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_19 <= io_in_weight_x_19; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_20 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_20 <= io_in_weight_x_20; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_21 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_21 <= io_in_weight_x_21; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_22 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_22 <= io_in_weight_x_22; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_23 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_23 <= io_in_weight_x_23; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_24 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_24 <= io_in_weight_x_24; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_25 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_25 <= io_in_weight_x_25; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_26 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_26 <= io_in_weight_x_26; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_27 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_27 <= io_in_weight_x_27; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_28 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_28 <= io_in_weight_x_28; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_29 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_29 <= io_in_weight_x_29; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_30 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_30 <= io_in_weight_x_30; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_31 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_31 <= io_in_weight_x_31; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_32 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_32 <= io_in_weight_x_32; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_33 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_33 <= io_in_weight_x_33; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_34 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_34 <= io_in_weight_x_34; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_35 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_35 <= io_in_weight_x_35; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_36 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_36 <= io_in_weight_x_36; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_37 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_37 <= io_in_weight_x_37; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_38 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_38 <= io_in_weight_x_38; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_39 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_39 <= io_in_weight_x_39; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_40 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_40 <= io_in_weight_x_40; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_41 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_41 <= io_in_weight_x_41; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_42 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_42 <= io_in_weight_x_42; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_43 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_43 <= io_in_weight_x_43; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_44 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_44 <= io_in_weight_x_44; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_45 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_45 <= io_in_weight_x_45; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_46 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_46 <= io_in_weight_x_46; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_47 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_47 <= io_in_weight_x_47; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_48 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_48 <= io_in_weight_x_48; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_49 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_49 <= io_in_weight_x_49; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_50 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_50 <= io_in_weight_x_50; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_51 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_51 <= io_in_weight_x_51; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_52 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_52 <= io_in_weight_x_52; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_53 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_53 <= io_in_weight_x_53; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_54 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_54 <= io_in_weight_x_54; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_55 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_55 <= io_in_weight_x_55; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_56 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_56 <= io_in_weight_x_56; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_57 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_57 <= io_in_weight_x_57; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_58 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_58 <= io_in_weight_x_58; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_59 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_59 <= io_in_weight_x_59; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_60 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_60 <= io_in_weight_x_60; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_61 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_61 <= io_in_weight_x_61; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_62 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_62 <= io_in_weight_x_62; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_1_63 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h1 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_1_63 <= io_in_weight_x_63; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_0 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_0 <= io_in_weight_x_0; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_1 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_1 <= io_in_weight_x_1; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_2 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_2 <= io_in_weight_x_2; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_3 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_3 <= io_in_weight_x_3; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_4 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_4 <= io_in_weight_x_4; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_5 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_5 <= io_in_weight_x_5; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_6 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_6 <= io_in_weight_x_6; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_7 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_7 <= io_in_weight_x_7; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_8 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_8 <= io_in_weight_x_8; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_9 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_9 <= io_in_weight_x_9; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_10 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_10 <= io_in_weight_x_10; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_11 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_11 <= io_in_weight_x_11; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_12 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_12 <= io_in_weight_x_12; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_13 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_13 <= io_in_weight_x_13; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_14 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_14 <= io_in_weight_x_14; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_15 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_15 <= io_in_weight_x_15; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_16 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_16 <= io_in_weight_x_16; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_17 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_17 <= io_in_weight_x_17; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_18 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_18 <= io_in_weight_x_18; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_19 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_19 <= io_in_weight_x_19; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_20 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_20 <= io_in_weight_x_20; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_21 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_21 <= io_in_weight_x_21; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_22 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_22 <= io_in_weight_x_22; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_23 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_23 <= io_in_weight_x_23; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_24 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_24 <= io_in_weight_x_24; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_25 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_25 <= io_in_weight_x_25; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_26 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_26 <= io_in_weight_x_26; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_27 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_27 <= io_in_weight_x_27; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_28 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_28 <= io_in_weight_x_28; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_29 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_29 <= io_in_weight_x_29; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_30 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_30 <= io_in_weight_x_30; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_31 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_31 <= io_in_weight_x_31; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_32 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_32 <= io_in_weight_x_32; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_33 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_33 <= io_in_weight_x_33; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_34 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_34 <= io_in_weight_x_34; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_35 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_35 <= io_in_weight_x_35; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_36 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_36 <= io_in_weight_x_36; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_37 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_37 <= io_in_weight_x_37; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_38 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_38 <= io_in_weight_x_38; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_39 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_39 <= io_in_weight_x_39; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_40 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_40 <= io_in_weight_x_40; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_41 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_41 <= io_in_weight_x_41; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_42 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_42 <= io_in_weight_x_42; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_43 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_43 <= io_in_weight_x_43; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_44 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_44 <= io_in_weight_x_44; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_45 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_45 <= io_in_weight_x_45; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_46 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_46 <= io_in_weight_x_46; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_47 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_47 <= io_in_weight_x_47; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_48 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_48 <= io_in_weight_x_48; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_49 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_49 <= io_in_weight_x_49; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_50 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_50 <= io_in_weight_x_50; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_51 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_51 <= io_in_weight_x_51; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_52 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_52 <= io_in_weight_x_52; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_53 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_53 <= io_in_weight_x_53; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_54 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_54 <= io_in_weight_x_54; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_55 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_55 <= io_in_weight_x_55; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_56 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_56 <= io_in_weight_x_56; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_57 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_57 <= io_in_weight_x_57; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_58 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_58 <= io_in_weight_x_58; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_59 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_59 <= io_in_weight_x_59; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_60 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_60 <= io_in_weight_x_60; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_61 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_61 <= io_in_weight_x_61; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_62 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_62 <= io_in_weight_x_62; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_2_63 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h2 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_2_63 <= io_in_weight_x_63; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_0 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_0 <= io_in_weight_x_0; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_1 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_1 <= io_in_weight_x_1; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_2 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_2 <= io_in_weight_x_2; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_3 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_3 <= io_in_weight_x_3; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_4 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_4 <= io_in_weight_x_4; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_5 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_5 <= io_in_weight_x_5; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_6 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_6 <= io_in_weight_x_6; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_7 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_7 <= io_in_weight_x_7; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_8 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_8 <= io_in_weight_x_8; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_9 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_9 <= io_in_weight_x_9; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_10 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_10 <= io_in_weight_x_10; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_11 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_11 <= io_in_weight_x_11; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_12 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_12 <= io_in_weight_x_12; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_13 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_13 <= io_in_weight_x_13; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_14 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_14 <= io_in_weight_x_14; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_15 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_15 <= io_in_weight_x_15; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_16 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_16 <= io_in_weight_x_16; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_17 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_17 <= io_in_weight_x_17; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_18 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_18 <= io_in_weight_x_18; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_19 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_19 <= io_in_weight_x_19; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_20 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_20 <= io_in_weight_x_20; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_21 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_21 <= io_in_weight_x_21; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_22 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_22 <= io_in_weight_x_22; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_23 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_23 <= io_in_weight_x_23; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_24 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_24 <= io_in_weight_x_24; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_25 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_25 <= io_in_weight_x_25; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_26 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_26 <= io_in_weight_x_26; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_27 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_27 <= io_in_weight_x_27; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_28 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_28 <= io_in_weight_x_28; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_29 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_29 <= io_in_weight_x_29; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_30 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_30 <= io_in_weight_x_30; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_31 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_31 <= io_in_weight_x_31; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_32 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_32 <= io_in_weight_x_32; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_33 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_33 <= io_in_weight_x_33; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_34 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_34 <= io_in_weight_x_34; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_35 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_35 <= io_in_weight_x_35; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_36 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_36 <= io_in_weight_x_36; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_37 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_37 <= io_in_weight_x_37; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_38 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_38 <= io_in_weight_x_38; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_39 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_39 <= io_in_weight_x_39; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_40 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_40 <= io_in_weight_x_40; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_41 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_41 <= io_in_weight_x_41; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_42 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_42 <= io_in_weight_x_42; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_43 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_43 <= io_in_weight_x_43; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_44 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_44 <= io_in_weight_x_44; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_45 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_45 <= io_in_weight_x_45; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_46 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_46 <= io_in_weight_x_46; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_47 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_47 <= io_in_weight_x_47; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_48 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_48 <= io_in_weight_x_48; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_49 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_49 <= io_in_weight_x_49; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_50 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_50 <= io_in_weight_x_50; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_51 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_51 <= io_in_weight_x_51; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_52 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_52 <= io_in_weight_x_52; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_53 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_53 <= io_in_weight_x_53; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_54 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_54 <= io_in_weight_x_54; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_55 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_55 <= io_in_weight_x_55; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_56 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_56 <= io_in_weight_x_56; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_57 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_57 <= io_in_weight_x_57; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_58 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_58 <= io_in_weight_x_58; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_59 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_59 <= io_in_weight_x_59; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_60 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_60 <= io_in_weight_x_60; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_61 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_61 <= io_in_weight_x_61; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_62 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_62 <= io_in_weight_x_62; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 25:23]
      buffer_3_63 <= 8'h0; // @[Weight_Buffer.scala 25:23]
    end else if (_T_1) begin // @[Weight_Buffer.scala 46:27]
      if (2'h3 == write_ptr[1:0]) begin // @[Weight_Buffer.scala 47:44]
        buffer_3_63 <= io_in_weight_x_63; // @[Weight_Buffer.scala 47:44]
      end
    end
    if (reset) begin // @[Weight_Buffer.scala 28:25]
      read_ptr <= 3'h0; // @[Weight_Buffer.scala 28:25]
    end else if (shift_ptr == 4'h0) begin // @[Weight_Buffer.scala 73:27]
      read_ptr <= _read_ptr_T_1; // @[Weight_Buffer.scala 74:14]
    end
    if (reset) begin // @[Weight_Buffer.scala 29:26]
      write_ptr <= 3'h0; // @[Weight_Buffer.scala 29:26]
    end else if (io_wen & ~full) begin // @[Weight_Buffer.scala 40:27]
      write_ptr <= _write_ptr_T_1; // @[Weight_Buffer.scala 41:15]
    end
    if (reset) begin // @[Weight_Buffer.scala 51:26]
      shift_ptr <= 4'h8; // @[Weight_Buffer.scala 51:26]
    end else if (io_ren & ~empty) begin // @[Weight_Buffer.scala 53:28]
      shift_ptr <= _shift_ptr_T_1; // @[Weight_Buffer.scala 54:15]
    end else if (4'h1 <= shift_ptr & shift_ptr < 4'h8) begin // @[Weight_Buffer.scala 55:61]
      shift_ptr <= _shift_ptr_T_1; // @[Weight_Buffer.scala 56:15]
    end else begin
      shift_ptr <= 4'h8; // @[Weight_Buffer.scala 58:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buffer_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_0_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_0_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_0_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_0_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_0_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_0_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_0_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_0_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_0_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_0_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_0_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_0_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_0_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_0_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_0_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_0_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_0_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_0_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_0_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_0_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_0_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_0_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_0_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_0_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_0_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_0_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_0_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_0_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_0_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_0_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_0_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_0_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_0_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_0_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_0_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_0_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_0_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_0_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_0_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_0_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_0_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_0_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_0_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_0_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  buffer_0_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_0_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_0_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_0_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_0_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  buffer_0_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_0_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_0_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_0_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_0_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  buffer_0_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_0_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_0_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_0_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_0_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  buffer_1_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_1_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_1_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_1_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_1_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  buffer_1_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_1_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_1_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_1_8 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_1_9 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  buffer_1_10 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_1_11 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_1_12 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_1_13 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  buffer_1_14 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  buffer_1_15 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_1_16 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_1_17 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  buffer_1_18 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  buffer_1_19 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  buffer_1_20 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  buffer_1_21 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  buffer_1_22 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  buffer_1_23 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  buffer_1_24 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  buffer_1_25 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  buffer_1_26 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  buffer_1_27 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  buffer_1_28 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  buffer_1_29 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  buffer_1_30 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  buffer_1_31 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  buffer_1_32 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  buffer_1_33 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  buffer_1_34 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  buffer_1_35 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  buffer_1_36 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  buffer_1_37 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  buffer_1_38 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  buffer_1_39 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  buffer_1_40 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  buffer_1_41 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  buffer_1_42 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  buffer_1_43 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  buffer_1_44 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  buffer_1_45 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  buffer_1_46 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  buffer_1_47 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  buffer_1_48 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  buffer_1_49 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  buffer_1_50 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  buffer_1_51 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  buffer_1_52 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  buffer_1_53 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  buffer_1_54 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  buffer_1_55 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  buffer_1_56 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  buffer_1_57 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  buffer_1_58 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  buffer_1_59 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  buffer_1_60 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  buffer_1_61 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  buffer_1_62 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  buffer_1_63 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  buffer_2_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  buffer_2_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  buffer_2_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  buffer_2_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  buffer_2_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  buffer_2_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  buffer_2_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  buffer_2_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  buffer_2_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  buffer_2_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  buffer_2_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  buffer_2_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  buffer_2_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  buffer_2_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  buffer_2_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  buffer_2_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  buffer_2_16 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  buffer_2_17 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  buffer_2_18 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  buffer_2_19 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  buffer_2_20 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  buffer_2_21 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  buffer_2_22 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  buffer_2_23 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  buffer_2_24 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  buffer_2_25 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  buffer_2_26 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  buffer_2_27 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  buffer_2_28 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  buffer_2_29 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  buffer_2_30 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  buffer_2_31 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  buffer_2_32 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  buffer_2_33 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  buffer_2_34 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  buffer_2_35 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  buffer_2_36 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  buffer_2_37 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  buffer_2_38 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  buffer_2_39 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  buffer_2_40 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  buffer_2_41 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  buffer_2_42 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  buffer_2_43 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  buffer_2_44 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  buffer_2_45 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  buffer_2_46 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  buffer_2_47 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  buffer_2_48 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  buffer_2_49 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  buffer_2_50 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  buffer_2_51 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  buffer_2_52 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  buffer_2_53 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  buffer_2_54 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  buffer_2_55 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  buffer_2_56 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  buffer_2_57 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  buffer_2_58 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  buffer_2_59 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  buffer_2_60 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  buffer_2_61 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  buffer_2_62 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  buffer_2_63 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  buffer_3_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  buffer_3_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  buffer_3_2 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  buffer_3_3 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  buffer_3_4 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  buffer_3_5 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  buffer_3_6 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  buffer_3_7 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  buffer_3_8 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  buffer_3_9 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  buffer_3_10 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  buffer_3_11 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  buffer_3_12 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  buffer_3_13 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  buffer_3_14 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  buffer_3_15 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  buffer_3_16 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  buffer_3_17 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  buffer_3_18 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  buffer_3_19 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  buffer_3_20 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  buffer_3_21 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  buffer_3_22 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  buffer_3_23 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  buffer_3_24 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  buffer_3_25 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  buffer_3_26 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  buffer_3_27 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  buffer_3_28 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  buffer_3_29 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  buffer_3_30 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  buffer_3_31 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  buffer_3_32 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  buffer_3_33 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  buffer_3_34 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  buffer_3_35 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  buffer_3_36 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  buffer_3_37 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  buffer_3_38 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  buffer_3_39 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  buffer_3_40 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  buffer_3_41 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  buffer_3_42 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  buffer_3_43 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  buffer_3_44 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  buffer_3_45 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  buffer_3_46 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  buffer_3_47 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  buffer_3_48 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  buffer_3_49 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  buffer_3_50 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  buffer_3_51 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  buffer_3_52 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  buffer_3_53 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  buffer_3_54 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  buffer_3_55 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  buffer_3_56 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  buffer_3_57 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  buffer_3_58 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  buffer_3_59 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  buffer_3_60 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  buffer_3_61 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  buffer_3_62 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  buffer_3_63 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  read_ptr = _RAND_256[2:0];
  _RAND_257 = {1{`RANDOM}};
  write_ptr = _RAND_257[2:0];
  _RAND_258 = {1{`RANDOM}};
  shift_ptr = _RAND_258[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module basic_PE(
  input         clock,
  input         reset,
  input  [7:0]  io_in_activate,
  input  [7:0]  io_in_weight,
  input  [15:0] io_in_psum,
  input         io_in_flow,
  input         io_in_shift,
  output [7:0]  io_out_activate,
  output [7:0]  io_out_weight,
  output [15:0] io_out_psum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] Activation_Reg; // @[basic_PE.scala 17:31]
  reg [7:0] Weight_Reg; // @[basic_PE.scala 18:27]
  reg [15:0] PSum_Reg; // @[basic_PE.scala 19:25]
  wire [15:0] _io_out_psum_T = Activation_Reg * Weight_Reg; // @[basic_PE.scala 47:33]
  assign io_out_activate = Activation_Reg; // @[basic_PE.scala 45:19]
  assign io_out_weight = Weight_Reg; // @[basic_PE.scala 46:17]
  assign io_out_psum = _io_out_psum_T + PSum_Reg; // @[basic_PE.scala 47:46]
  always @(posedge clock) begin
    if (reset) begin // @[basic_PE.scala 17:31]
      Activation_Reg <= 8'h0; // @[basic_PE.scala 17:31]
    end else if (io_in_flow) begin // @[basic_PE.scala 22:20]
      Activation_Reg <= io_in_activate; // @[basic_PE.scala 23:20]
    end
    if (reset) begin // @[basic_PE.scala 18:27]
      Weight_Reg <= 8'h0; // @[basic_PE.scala 18:27]
    end else if (io_in_shift) begin // @[basic_PE.scala 38:21]
      Weight_Reg <= io_in_weight; // @[basic_PE.scala 39:16]
    end
    if (reset) begin // @[basic_PE.scala 19:25]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 19:25]
    end else if (io_in_shift) begin // @[basic_PE.scala 29:21]
      PSum_Reg <= 16'h0; // @[basic_PE.scala 30:14]
    end else if (io_in_flow) begin // @[basic_PE.scala 31:26]
      PSum_Reg <= io_in_psum; // @[basic_PE.scala 32:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Activation_Reg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  Weight_Reg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  PSum_Reg = _RAND_2[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Systolic_Array(
  input         clock,
  input         reset,
  input  [7:0]  io_activate_0,
  input  [7:0]  io_activate_1,
  input  [7:0]  io_activate_2,
  input  [7:0]  io_activate_3,
  input  [7:0]  io_activate_4,
  input  [7:0]  io_activate_5,
  input  [7:0]  io_activate_6,
  input  [7:0]  io_activate_7,
  input  [7:0]  io_weight_0,
  input  [7:0]  io_weight_1,
  input  [7:0]  io_weight_2,
  input  [7:0]  io_weight_3,
  input  [7:0]  io_weight_4,
  input  [7:0]  io_weight_5,
  input  [7:0]  io_weight_6,
  input  [7:0]  io_weight_7,
  input         io_flow,
  input         io_shift,
  output [15:0] io_psum_0,
  output [15:0] io_psum_1,
  output [15:0] io_psum_2,
  output [15:0] io_psum_3,
  output [15:0] io_psum_4,
  output [15:0] io_psum_5,
  output [15:0] io_psum_6,
  output [15:0] io_psum_7,
  output        io_valid_0,
  output        io_valid_1,
  output        io_valid_2,
  output        io_valid_3,
  output        io_valid_4,
  output        io_valid_5,
  output        io_valid_6,
  output        io_valid_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  PE_Array_0_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_0_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_0_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_0_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_1_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_1_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_1_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_2_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_2_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_2_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_3_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_3_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_3_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_4_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_4_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_4_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_5_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_5_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_5_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_6_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_6_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_6_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_0_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_0_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_0_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_1_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_1_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_1_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_2_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_2_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_2_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_3_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_3_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_3_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_4_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_4_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_4_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_5_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_5_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_5_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_6_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_6_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_6_io_out_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_clock; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_reset; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_in_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_in_psum; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_flow; // @[Systolic_Array.scala 19:62]
  wire  PE_Array_7_7_io_in_shift; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_activate; // @[Systolic_Array.scala 19:62]
  wire [7:0] PE_Array_7_7_io_out_weight; // @[Systolic_Array.scala 19:62]
  wire [15:0] PE_Array_7_7_io_out_psum; // @[Systolic_Array.scala 19:62]
  reg [4:0] flow_counter; // @[Systolic_Array.scala 52:29]
  reg [7:0] valid_reg; // @[Systolic_Array.scala 53:26]
  wire [4:0] _flow_counter_T_1 = flow_counter + 5'h1; // @[Systolic_Array.scala 57:34]
  wire [7:0] _valid_reg_T_1 = {valid_reg[6:0],1'h1}; // @[Cat.scala 33:92]
  wire [7:0] _valid_reg_T_3 = {valid_reg[6:0],1'h0}; // @[Cat.scala 33:92]
  basic_PE PE_Array_0_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_0_clock),
    .reset(PE_Array_0_0_reset),
    .io_in_activate(PE_Array_0_0_io_in_activate),
    .io_in_weight(PE_Array_0_0_io_in_weight),
    .io_in_psum(PE_Array_0_0_io_in_psum),
    .io_in_flow(PE_Array_0_0_io_in_flow),
    .io_in_shift(PE_Array_0_0_io_in_shift),
    .io_out_activate(PE_Array_0_0_io_out_activate),
    .io_out_weight(PE_Array_0_0_io_out_weight),
    .io_out_psum(PE_Array_0_0_io_out_psum)
  );
  basic_PE PE_Array_0_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_1_clock),
    .reset(PE_Array_0_1_reset),
    .io_in_activate(PE_Array_0_1_io_in_activate),
    .io_in_weight(PE_Array_0_1_io_in_weight),
    .io_in_psum(PE_Array_0_1_io_in_psum),
    .io_in_flow(PE_Array_0_1_io_in_flow),
    .io_in_shift(PE_Array_0_1_io_in_shift),
    .io_out_activate(PE_Array_0_1_io_out_activate),
    .io_out_weight(PE_Array_0_1_io_out_weight),
    .io_out_psum(PE_Array_0_1_io_out_psum)
  );
  basic_PE PE_Array_0_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_2_clock),
    .reset(PE_Array_0_2_reset),
    .io_in_activate(PE_Array_0_2_io_in_activate),
    .io_in_weight(PE_Array_0_2_io_in_weight),
    .io_in_psum(PE_Array_0_2_io_in_psum),
    .io_in_flow(PE_Array_0_2_io_in_flow),
    .io_in_shift(PE_Array_0_2_io_in_shift),
    .io_out_activate(PE_Array_0_2_io_out_activate),
    .io_out_weight(PE_Array_0_2_io_out_weight),
    .io_out_psum(PE_Array_0_2_io_out_psum)
  );
  basic_PE PE_Array_0_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_3_clock),
    .reset(PE_Array_0_3_reset),
    .io_in_activate(PE_Array_0_3_io_in_activate),
    .io_in_weight(PE_Array_0_3_io_in_weight),
    .io_in_psum(PE_Array_0_3_io_in_psum),
    .io_in_flow(PE_Array_0_3_io_in_flow),
    .io_in_shift(PE_Array_0_3_io_in_shift),
    .io_out_activate(PE_Array_0_3_io_out_activate),
    .io_out_weight(PE_Array_0_3_io_out_weight),
    .io_out_psum(PE_Array_0_3_io_out_psum)
  );
  basic_PE PE_Array_0_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_4_clock),
    .reset(PE_Array_0_4_reset),
    .io_in_activate(PE_Array_0_4_io_in_activate),
    .io_in_weight(PE_Array_0_4_io_in_weight),
    .io_in_psum(PE_Array_0_4_io_in_psum),
    .io_in_flow(PE_Array_0_4_io_in_flow),
    .io_in_shift(PE_Array_0_4_io_in_shift),
    .io_out_activate(PE_Array_0_4_io_out_activate),
    .io_out_weight(PE_Array_0_4_io_out_weight),
    .io_out_psum(PE_Array_0_4_io_out_psum)
  );
  basic_PE PE_Array_0_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_5_clock),
    .reset(PE_Array_0_5_reset),
    .io_in_activate(PE_Array_0_5_io_in_activate),
    .io_in_weight(PE_Array_0_5_io_in_weight),
    .io_in_psum(PE_Array_0_5_io_in_psum),
    .io_in_flow(PE_Array_0_5_io_in_flow),
    .io_in_shift(PE_Array_0_5_io_in_shift),
    .io_out_activate(PE_Array_0_5_io_out_activate),
    .io_out_weight(PE_Array_0_5_io_out_weight),
    .io_out_psum(PE_Array_0_5_io_out_psum)
  );
  basic_PE PE_Array_0_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_6_clock),
    .reset(PE_Array_0_6_reset),
    .io_in_activate(PE_Array_0_6_io_in_activate),
    .io_in_weight(PE_Array_0_6_io_in_weight),
    .io_in_psum(PE_Array_0_6_io_in_psum),
    .io_in_flow(PE_Array_0_6_io_in_flow),
    .io_in_shift(PE_Array_0_6_io_in_shift),
    .io_out_activate(PE_Array_0_6_io_out_activate),
    .io_out_weight(PE_Array_0_6_io_out_weight),
    .io_out_psum(PE_Array_0_6_io_out_psum)
  );
  basic_PE PE_Array_0_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_0_7_clock),
    .reset(PE_Array_0_7_reset),
    .io_in_activate(PE_Array_0_7_io_in_activate),
    .io_in_weight(PE_Array_0_7_io_in_weight),
    .io_in_psum(PE_Array_0_7_io_in_psum),
    .io_in_flow(PE_Array_0_7_io_in_flow),
    .io_in_shift(PE_Array_0_7_io_in_shift),
    .io_out_activate(PE_Array_0_7_io_out_activate),
    .io_out_weight(PE_Array_0_7_io_out_weight),
    .io_out_psum(PE_Array_0_7_io_out_psum)
  );
  basic_PE PE_Array_1_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_0_clock),
    .reset(PE_Array_1_0_reset),
    .io_in_activate(PE_Array_1_0_io_in_activate),
    .io_in_weight(PE_Array_1_0_io_in_weight),
    .io_in_psum(PE_Array_1_0_io_in_psum),
    .io_in_flow(PE_Array_1_0_io_in_flow),
    .io_in_shift(PE_Array_1_0_io_in_shift),
    .io_out_activate(PE_Array_1_0_io_out_activate),
    .io_out_weight(PE_Array_1_0_io_out_weight),
    .io_out_psum(PE_Array_1_0_io_out_psum)
  );
  basic_PE PE_Array_1_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_1_clock),
    .reset(PE_Array_1_1_reset),
    .io_in_activate(PE_Array_1_1_io_in_activate),
    .io_in_weight(PE_Array_1_1_io_in_weight),
    .io_in_psum(PE_Array_1_1_io_in_psum),
    .io_in_flow(PE_Array_1_1_io_in_flow),
    .io_in_shift(PE_Array_1_1_io_in_shift),
    .io_out_activate(PE_Array_1_1_io_out_activate),
    .io_out_weight(PE_Array_1_1_io_out_weight),
    .io_out_psum(PE_Array_1_1_io_out_psum)
  );
  basic_PE PE_Array_1_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_2_clock),
    .reset(PE_Array_1_2_reset),
    .io_in_activate(PE_Array_1_2_io_in_activate),
    .io_in_weight(PE_Array_1_2_io_in_weight),
    .io_in_psum(PE_Array_1_2_io_in_psum),
    .io_in_flow(PE_Array_1_2_io_in_flow),
    .io_in_shift(PE_Array_1_2_io_in_shift),
    .io_out_activate(PE_Array_1_2_io_out_activate),
    .io_out_weight(PE_Array_1_2_io_out_weight),
    .io_out_psum(PE_Array_1_2_io_out_psum)
  );
  basic_PE PE_Array_1_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_3_clock),
    .reset(PE_Array_1_3_reset),
    .io_in_activate(PE_Array_1_3_io_in_activate),
    .io_in_weight(PE_Array_1_3_io_in_weight),
    .io_in_psum(PE_Array_1_3_io_in_psum),
    .io_in_flow(PE_Array_1_3_io_in_flow),
    .io_in_shift(PE_Array_1_3_io_in_shift),
    .io_out_activate(PE_Array_1_3_io_out_activate),
    .io_out_weight(PE_Array_1_3_io_out_weight),
    .io_out_psum(PE_Array_1_3_io_out_psum)
  );
  basic_PE PE_Array_1_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_4_clock),
    .reset(PE_Array_1_4_reset),
    .io_in_activate(PE_Array_1_4_io_in_activate),
    .io_in_weight(PE_Array_1_4_io_in_weight),
    .io_in_psum(PE_Array_1_4_io_in_psum),
    .io_in_flow(PE_Array_1_4_io_in_flow),
    .io_in_shift(PE_Array_1_4_io_in_shift),
    .io_out_activate(PE_Array_1_4_io_out_activate),
    .io_out_weight(PE_Array_1_4_io_out_weight),
    .io_out_psum(PE_Array_1_4_io_out_psum)
  );
  basic_PE PE_Array_1_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_5_clock),
    .reset(PE_Array_1_5_reset),
    .io_in_activate(PE_Array_1_5_io_in_activate),
    .io_in_weight(PE_Array_1_5_io_in_weight),
    .io_in_psum(PE_Array_1_5_io_in_psum),
    .io_in_flow(PE_Array_1_5_io_in_flow),
    .io_in_shift(PE_Array_1_5_io_in_shift),
    .io_out_activate(PE_Array_1_5_io_out_activate),
    .io_out_weight(PE_Array_1_5_io_out_weight),
    .io_out_psum(PE_Array_1_5_io_out_psum)
  );
  basic_PE PE_Array_1_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_6_clock),
    .reset(PE_Array_1_6_reset),
    .io_in_activate(PE_Array_1_6_io_in_activate),
    .io_in_weight(PE_Array_1_6_io_in_weight),
    .io_in_psum(PE_Array_1_6_io_in_psum),
    .io_in_flow(PE_Array_1_6_io_in_flow),
    .io_in_shift(PE_Array_1_6_io_in_shift),
    .io_out_activate(PE_Array_1_6_io_out_activate),
    .io_out_weight(PE_Array_1_6_io_out_weight),
    .io_out_psum(PE_Array_1_6_io_out_psum)
  );
  basic_PE PE_Array_1_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_1_7_clock),
    .reset(PE_Array_1_7_reset),
    .io_in_activate(PE_Array_1_7_io_in_activate),
    .io_in_weight(PE_Array_1_7_io_in_weight),
    .io_in_psum(PE_Array_1_7_io_in_psum),
    .io_in_flow(PE_Array_1_7_io_in_flow),
    .io_in_shift(PE_Array_1_7_io_in_shift),
    .io_out_activate(PE_Array_1_7_io_out_activate),
    .io_out_weight(PE_Array_1_7_io_out_weight),
    .io_out_psum(PE_Array_1_7_io_out_psum)
  );
  basic_PE PE_Array_2_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_0_clock),
    .reset(PE_Array_2_0_reset),
    .io_in_activate(PE_Array_2_0_io_in_activate),
    .io_in_weight(PE_Array_2_0_io_in_weight),
    .io_in_psum(PE_Array_2_0_io_in_psum),
    .io_in_flow(PE_Array_2_0_io_in_flow),
    .io_in_shift(PE_Array_2_0_io_in_shift),
    .io_out_activate(PE_Array_2_0_io_out_activate),
    .io_out_weight(PE_Array_2_0_io_out_weight),
    .io_out_psum(PE_Array_2_0_io_out_psum)
  );
  basic_PE PE_Array_2_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_1_clock),
    .reset(PE_Array_2_1_reset),
    .io_in_activate(PE_Array_2_1_io_in_activate),
    .io_in_weight(PE_Array_2_1_io_in_weight),
    .io_in_psum(PE_Array_2_1_io_in_psum),
    .io_in_flow(PE_Array_2_1_io_in_flow),
    .io_in_shift(PE_Array_2_1_io_in_shift),
    .io_out_activate(PE_Array_2_1_io_out_activate),
    .io_out_weight(PE_Array_2_1_io_out_weight),
    .io_out_psum(PE_Array_2_1_io_out_psum)
  );
  basic_PE PE_Array_2_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_2_clock),
    .reset(PE_Array_2_2_reset),
    .io_in_activate(PE_Array_2_2_io_in_activate),
    .io_in_weight(PE_Array_2_2_io_in_weight),
    .io_in_psum(PE_Array_2_2_io_in_psum),
    .io_in_flow(PE_Array_2_2_io_in_flow),
    .io_in_shift(PE_Array_2_2_io_in_shift),
    .io_out_activate(PE_Array_2_2_io_out_activate),
    .io_out_weight(PE_Array_2_2_io_out_weight),
    .io_out_psum(PE_Array_2_2_io_out_psum)
  );
  basic_PE PE_Array_2_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_3_clock),
    .reset(PE_Array_2_3_reset),
    .io_in_activate(PE_Array_2_3_io_in_activate),
    .io_in_weight(PE_Array_2_3_io_in_weight),
    .io_in_psum(PE_Array_2_3_io_in_psum),
    .io_in_flow(PE_Array_2_3_io_in_flow),
    .io_in_shift(PE_Array_2_3_io_in_shift),
    .io_out_activate(PE_Array_2_3_io_out_activate),
    .io_out_weight(PE_Array_2_3_io_out_weight),
    .io_out_psum(PE_Array_2_3_io_out_psum)
  );
  basic_PE PE_Array_2_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_4_clock),
    .reset(PE_Array_2_4_reset),
    .io_in_activate(PE_Array_2_4_io_in_activate),
    .io_in_weight(PE_Array_2_4_io_in_weight),
    .io_in_psum(PE_Array_2_4_io_in_psum),
    .io_in_flow(PE_Array_2_4_io_in_flow),
    .io_in_shift(PE_Array_2_4_io_in_shift),
    .io_out_activate(PE_Array_2_4_io_out_activate),
    .io_out_weight(PE_Array_2_4_io_out_weight),
    .io_out_psum(PE_Array_2_4_io_out_psum)
  );
  basic_PE PE_Array_2_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_5_clock),
    .reset(PE_Array_2_5_reset),
    .io_in_activate(PE_Array_2_5_io_in_activate),
    .io_in_weight(PE_Array_2_5_io_in_weight),
    .io_in_psum(PE_Array_2_5_io_in_psum),
    .io_in_flow(PE_Array_2_5_io_in_flow),
    .io_in_shift(PE_Array_2_5_io_in_shift),
    .io_out_activate(PE_Array_2_5_io_out_activate),
    .io_out_weight(PE_Array_2_5_io_out_weight),
    .io_out_psum(PE_Array_2_5_io_out_psum)
  );
  basic_PE PE_Array_2_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_6_clock),
    .reset(PE_Array_2_6_reset),
    .io_in_activate(PE_Array_2_6_io_in_activate),
    .io_in_weight(PE_Array_2_6_io_in_weight),
    .io_in_psum(PE_Array_2_6_io_in_psum),
    .io_in_flow(PE_Array_2_6_io_in_flow),
    .io_in_shift(PE_Array_2_6_io_in_shift),
    .io_out_activate(PE_Array_2_6_io_out_activate),
    .io_out_weight(PE_Array_2_6_io_out_weight),
    .io_out_psum(PE_Array_2_6_io_out_psum)
  );
  basic_PE PE_Array_2_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_2_7_clock),
    .reset(PE_Array_2_7_reset),
    .io_in_activate(PE_Array_2_7_io_in_activate),
    .io_in_weight(PE_Array_2_7_io_in_weight),
    .io_in_psum(PE_Array_2_7_io_in_psum),
    .io_in_flow(PE_Array_2_7_io_in_flow),
    .io_in_shift(PE_Array_2_7_io_in_shift),
    .io_out_activate(PE_Array_2_7_io_out_activate),
    .io_out_weight(PE_Array_2_7_io_out_weight),
    .io_out_psum(PE_Array_2_7_io_out_psum)
  );
  basic_PE PE_Array_3_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_0_clock),
    .reset(PE_Array_3_0_reset),
    .io_in_activate(PE_Array_3_0_io_in_activate),
    .io_in_weight(PE_Array_3_0_io_in_weight),
    .io_in_psum(PE_Array_3_0_io_in_psum),
    .io_in_flow(PE_Array_3_0_io_in_flow),
    .io_in_shift(PE_Array_3_0_io_in_shift),
    .io_out_activate(PE_Array_3_0_io_out_activate),
    .io_out_weight(PE_Array_3_0_io_out_weight),
    .io_out_psum(PE_Array_3_0_io_out_psum)
  );
  basic_PE PE_Array_3_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_1_clock),
    .reset(PE_Array_3_1_reset),
    .io_in_activate(PE_Array_3_1_io_in_activate),
    .io_in_weight(PE_Array_3_1_io_in_weight),
    .io_in_psum(PE_Array_3_1_io_in_psum),
    .io_in_flow(PE_Array_3_1_io_in_flow),
    .io_in_shift(PE_Array_3_1_io_in_shift),
    .io_out_activate(PE_Array_3_1_io_out_activate),
    .io_out_weight(PE_Array_3_1_io_out_weight),
    .io_out_psum(PE_Array_3_1_io_out_psum)
  );
  basic_PE PE_Array_3_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_2_clock),
    .reset(PE_Array_3_2_reset),
    .io_in_activate(PE_Array_3_2_io_in_activate),
    .io_in_weight(PE_Array_3_2_io_in_weight),
    .io_in_psum(PE_Array_3_2_io_in_psum),
    .io_in_flow(PE_Array_3_2_io_in_flow),
    .io_in_shift(PE_Array_3_2_io_in_shift),
    .io_out_activate(PE_Array_3_2_io_out_activate),
    .io_out_weight(PE_Array_3_2_io_out_weight),
    .io_out_psum(PE_Array_3_2_io_out_psum)
  );
  basic_PE PE_Array_3_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_3_clock),
    .reset(PE_Array_3_3_reset),
    .io_in_activate(PE_Array_3_3_io_in_activate),
    .io_in_weight(PE_Array_3_3_io_in_weight),
    .io_in_psum(PE_Array_3_3_io_in_psum),
    .io_in_flow(PE_Array_3_3_io_in_flow),
    .io_in_shift(PE_Array_3_3_io_in_shift),
    .io_out_activate(PE_Array_3_3_io_out_activate),
    .io_out_weight(PE_Array_3_3_io_out_weight),
    .io_out_psum(PE_Array_3_3_io_out_psum)
  );
  basic_PE PE_Array_3_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_4_clock),
    .reset(PE_Array_3_4_reset),
    .io_in_activate(PE_Array_3_4_io_in_activate),
    .io_in_weight(PE_Array_3_4_io_in_weight),
    .io_in_psum(PE_Array_3_4_io_in_psum),
    .io_in_flow(PE_Array_3_4_io_in_flow),
    .io_in_shift(PE_Array_3_4_io_in_shift),
    .io_out_activate(PE_Array_3_4_io_out_activate),
    .io_out_weight(PE_Array_3_4_io_out_weight),
    .io_out_psum(PE_Array_3_4_io_out_psum)
  );
  basic_PE PE_Array_3_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_5_clock),
    .reset(PE_Array_3_5_reset),
    .io_in_activate(PE_Array_3_5_io_in_activate),
    .io_in_weight(PE_Array_3_5_io_in_weight),
    .io_in_psum(PE_Array_3_5_io_in_psum),
    .io_in_flow(PE_Array_3_5_io_in_flow),
    .io_in_shift(PE_Array_3_5_io_in_shift),
    .io_out_activate(PE_Array_3_5_io_out_activate),
    .io_out_weight(PE_Array_3_5_io_out_weight),
    .io_out_psum(PE_Array_3_5_io_out_psum)
  );
  basic_PE PE_Array_3_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_6_clock),
    .reset(PE_Array_3_6_reset),
    .io_in_activate(PE_Array_3_6_io_in_activate),
    .io_in_weight(PE_Array_3_6_io_in_weight),
    .io_in_psum(PE_Array_3_6_io_in_psum),
    .io_in_flow(PE_Array_3_6_io_in_flow),
    .io_in_shift(PE_Array_3_6_io_in_shift),
    .io_out_activate(PE_Array_3_6_io_out_activate),
    .io_out_weight(PE_Array_3_6_io_out_weight),
    .io_out_psum(PE_Array_3_6_io_out_psum)
  );
  basic_PE PE_Array_3_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_3_7_clock),
    .reset(PE_Array_3_7_reset),
    .io_in_activate(PE_Array_3_7_io_in_activate),
    .io_in_weight(PE_Array_3_7_io_in_weight),
    .io_in_psum(PE_Array_3_7_io_in_psum),
    .io_in_flow(PE_Array_3_7_io_in_flow),
    .io_in_shift(PE_Array_3_7_io_in_shift),
    .io_out_activate(PE_Array_3_7_io_out_activate),
    .io_out_weight(PE_Array_3_7_io_out_weight),
    .io_out_psum(PE_Array_3_7_io_out_psum)
  );
  basic_PE PE_Array_4_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_0_clock),
    .reset(PE_Array_4_0_reset),
    .io_in_activate(PE_Array_4_0_io_in_activate),
    .io_in_weight(PE_Array_4_0_io_in_weight),
    .io_in_psum(PE_Array_4_0_io_in_psum),
    .io_in_flow(PE_Array_4_0_io_in_flow),
    .io_in_shift(PE_Array_4_0_io_in_shift),
    .io_out_activate(PE_Array_4_0_io_out_activate),
    .io_out_weight(PE_Array_4_0_io_out_weight),
    .io_out_psum(PE_Array_4_0_io_out_psum)
  );
  basic_PE PE_Array_4_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_1_clock),
    .reset(PE_Array_4_1_reset),
    .io_in_activate(PE_Array_4_1_io_in_activate),
    .io_in_weight(PE_Array_4_1_io_in_weight),
    .io_in_psum(PE_Array_4_1_io_in_psum),
    .io_in_flow(PE_Array_4_1_io_in_flow),
    .io_in_shift(PE_Array_4_1_io_in_shift),
    .io_out_activate(PE_Array_4_1_io_out_activate),
    .io_out_weight(PE_Array_4_1_io_out_weight),
    .io_out_psum(PE_Array_4_1_io_out_psum)
  );
  basic_PE PE_Array_4_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_2_clock),
    .reset(PE_Array_4_2_reset),
    .io_in_activate(PE_Array_4_2_io_in_activate),
    .io_in_weight(PE_Array_4_2_io_in_weight),
    .io_in_psum(PE_Array_4_2_io_in_psum),
    .io_in_flow(PE_Array_4_2_io_in_flow),
    .io_in_shift(PE_Array_4_2_io_in_shift),
    .io_out_activate(PE_Array_4_2_io_out_activate),
    .io_out_weight(PE_Array_4_2_io_out_weight),
    .io_out_psum(PE_Array_4_2_io_out_psum)
  );
  basic_PE PE_Array_4_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_3_clock),
    .reset(PE_Array_4_3_reset),
    .io_in_activate(PE_Array_4_3_io_in_activate),
    .io_in_weight(PE_Array_4_3_io_in_weight),
    .io_in_psum(PE_Array_4_3_io_in_psum),
    .io_in_flow(PE_Array_4_3_io_in_flow),
    .io_in_shift(PE_Array_4_3_io_in_shift),
    .io_out_activate(PE_Array_4_3_io_out_activate),
    .io_out_weight(PE_Array_4_3_io_out_weight),
    .io_out_psum(PE_Array_4_3_io_out_psum)
  );
  basic_PE PE_Array_4_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_4_clock),
    .reset(PE_Array_4_4_reset),
    .io_in_activate(PE_Array_4_4_io_in_activate),
    .io_in_weight(PE_Array_4_4_io_in_weight),
    .io_in_psum(PE_Array_4_4_io_in_psum),
    .io_in_flow(PE_Array_4_4_io_in_flow),
    .io_in_shift(PE_Array_4_4_io_in_shift),
    .io_out_activate(PE_Array_4_4_io_out_activate),
    .io_out_weight(PE_Array_4_4_io_out_weight),
    .io_out_psum(PE_Array_4_4_io_out_psum)
  );
  basic_PE PE_Array_4_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_5_clock),
    .reset(PE_Array_4_5_reset),
    .io_in_activate(PE_Array_4_5_io_in_activate),
    .io_in_weight(PE_Array_4_5_io_in_weight),
    .io_in_psum(PE_Array_4_5_io_in_psum),
    .io_in_flow(PE_Array_4_5_io_in_flow),
    .io_in_shift(PE_Array_4_5_io_in_shift),
    .io_out_activate(PE_Array_4_5_io_out_activate),
    .io_out_weight(PE_Array_4_5_io_out_weight),
    .io_out_psum(PE_Array_4_5_io_out_psum)
  );
  basic_PE PE_Array_4_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_6_clock),
    .reset(PE_Array_4_6_reset),
    .io_in_activate(PE_Array_4_6_io_in_activate),
    .io_in_weight(PE_Array_4_6_io_in_weight),
    .io_in_psum(PE_Array_4_6_io_in_psum),
    .io_in_flow(PE_Array_4_6_io_in_flow),
    .io_in_shift(PE_Array_4_6_io_in_shift),
    .io_out_activate(PE_Array_4_6_io_out_activate),
    .io_out_weight(PE_Array_4_6_io_out_weight),
    .io_out_psum(PE_Array_4_6_io_out_psum)
  );
  basic_PE PE_Array_4_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_4_7_clock),
    .reset(PE_Array_4_7_reset),
    .io_in_activate(PE_Array_4_7_io_in_activate),
    .io_in_weight(PE_Array_4_7_io_in_weight),
    .io_in_psum(PE_Array_4_7_io_in_psum),
    .io_in_flow(PE_Array_4_7_io_in_flow),
    .io_in_shift(PE_Array_4_7_io_in_shift),
    .io_out_activate(PE_Array_4_7_io_out_activate),
    .io_out_weight(PE_Array_4_7_io_out_weight),
    .io_out_psum(PE_Array_4_7_io_out_psum)
  );
  basic_PE PE_Array_5_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_0_clock),
    .reset(PE_Array_5_0_reset),
    .io_in_activate(PE_Array_5_0_io_in_activate),
    .io_in_weight(PE_Array_5_0_io_in_weight),
    .io_in_psum(PE_Array_5_0_io_in_psum),
    .io_in_flow(PE_Array_5_0_io_in_flow),
    .io_in_shift(PE_Array_5_0_io_in_shift),
    .io_out_activate(PE_Array_5_0_io_out_activate),
    .io_out_weight(PE_Array_5_0_io_out_weight),
    .io_out_psum(PE_Array_5_0_io_out_psum)
  );
  basic_PE PE_Array_5_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_1_clock),
    .reset(PE_Array_5_1_reset),
    .io_in_activate(PE_Array_5_1_io_in_activate),
    .io_in_weight(PE_Array_5_1_io_in_weight),
    .io_in_psum(PE_Array_5_1_io_in_psum),
    .io_in_flow(PE_Array_5_1_io_in_flow),
    .io_in_shift(PE_Array_5_1_io_in_shift),
    .io_out_activate(PE_Array_5_1_io_out_activate),
    .io_out_weight(PE_Array_5_1_io_out_weight),
    .io_out_psum(PE_Array_5_1_io_out_psum)
  );
  basic_PE PE_Array_5_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_2_clock),
    .reset(PE_Array_5_2_reset),
    .io_in_activate(PE_Array_5_2_io_in_activate),
    .io_in_weight(PE_Array_5_2_io_in_weight),
    .io_in_psum(PE_Array_5_2_io_in_psum),
    .io_in_flow(PE_Array_5_2_io_in_flow),
    .io_in_shift(PE_Array_5_2_io_in_shift),
    .io_out_activate(PE_Array_5_2_io_out_activate),
    .io_out_weight(PE_Array_5_2_io_out_weight),
    .io_out_psum(PE_Array_5_2_io_out_psum)
  );
  basic_PE PE_Array_5_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_3_clock),
    .reset(PE_Array_5_3_reset),
    .io_in_activate(PE_Array_5_3_io_in_activate),
    .io_in_weight(PE_Array_5_3_io_in_weight),
    .io_in_psum(PE_Array_5_3_io_in_psum),
    .io_in_flow(PE_Array_5_3_io_in_flow),
    .io_in_shift(PE_Array_5_3_io_in_shift),
    .io_out_activate(PE_Array_5_3_io_out_activate),
    .io_out_weight(PE_Array_5_3_io_out_weight),
    .io_out_psum(PE_Array_5_3_io_out_psum)
  );
  basic_PE PE_Array_5_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_4_clock),
    .reset(PE_Array_5_4_reset),
    .io_in_activate(PE_Array_5_4_io_in_activate),
    .io_in_weight(PE_Array_5_4_io_in_weight),
    .io_in_psum(PE_Array_5_4_io_in_psum),
    .io_in_flow(PE_Array_5_4_io_in_flow),
    .io_in_shift(PE_Array_5_4_io_in_shift),
    .io_out_activate(PE_Array_5_4_io_out_activate),
    .io_out_weight(PE_Array_5_4_io_out_weight),
    .io_out_psum(PE_Array_5_4_io_out_psum)
  );
  basic_PE PE_Array_5_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_5_clock),
    .reset(PE_Array_5_5_reset),
    .io_in_activate(PE_Array_5_5_io_in_activate),
    .io_in_weight(PE_Array_5_5_io_in_weight),
    .io_in_psum(PE_Array_5_5_io_in_psum),
    .io_in_flow(PE_Array_5_5_io_in_flow),
    .io_in_shift(PE_Array_5_5_io_in_shift),
    .io_out_activate(PE_Array_5_5_io_out_activate),
    .io_out_weight(PE_Array_5_5_io_out_weight),
    .io_out_psum(PE_Array_5_5_io_out_psum)
  );
  basic_PE PE_Array_5_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_6_clock),
    .reset(PE_Array_5_6_reset),
    .io_in_activate(PE_Array_5_6_io_in_activate),
    .io_in_weight(PE_Array_5_6_io_in_weight),
    .io_in_psum(PE_Array_5_6_io_in_psum),
    .io_in_flow(PE_Array_5_6_io_in_flow),
    .io_in_shift(PE_Array_5_6_io_in_shift),
    .io_out_activate(PE_Array_5_6_io_out_activate),
    .io_out_weight(PE_Array_5_6_io_out_weight),
    .io_out_psum(PE_Array_5_6_io_out_psum)
  );
  basic_PE PE_Array_5_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_5_7_clock),
    .reset(PE_Array_5_7_reset),
    .io_in_activate(PE_Array_5_7_io_in_activate),
    .io_in_weight(PE_Array_5_7_io_in_weight),
    .io_in_psum(PE_Array_5_7_io_in_psum),
    .io_in_flow(PE_Array_5_7_io_in_flow),
    .io_in_shift(PE_Array_5_7_io_in_shift),
    .io_out_activate(PE_Array_5_7_io_out_activate),
    .io_out_weight(PE_Array_5_7_io_out_weight),
    .io_out_psum(PE_Array_5_7_io_out_psum)
  );
  basic_PE PE_Array_6_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_0_clock),
    .reset(PE_Array_6_0_reset),
    .io_in_activate(PE_Array_6_0_io_in_activate),
    .io_in_weight(PE_Array_6_0_io_in_weight),
    .io_in_psum(PE_Array_6_0_io_in_psum),
    .io_in_flow(PE_Array_6_0_io_in_flow),
    .io_in_shift(PE_Array_6_0_io_in_shift),
    .io_out_activate(PE_Array_6_0_io_out_activate),
    .io_out_weight(PE_Array_6_0_io_out_weight),
    .io_out_psum(PE_Array_6_0_io_out_psum)
  );
  basic_PE PE_Array_6_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_1_clock),
    .reset(PE_Array_6_1_reset),
    .io_in_activate(PE_Array_6_1_io_in_activate),
    .io_in_weight(PE_Array_6_1_io_in_weight),
    .io_in_psum(PE_Array_6_1_io_in_psum),
    .io_in_flow(PE_Array_6_1_io_in_flow),
    .io_in_shift(PE_Array_6_1_io_in_shift),
    .io_out_activate(PE_Array_6_1_io_out_activate),
    .io_out_weight(PE_Array_6_1_io_out_weight),
    .io_out_psum(PE_Array_6_1_io_out_psum)
  );
  basic_PE PE_Array_6_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_2_clock),
    .reset(PE_Array_6_2_reset),
    .io_in_activate(PE_Array_6_2_io_in_activate),
    .io_in_weight(PE_Array_6_2_io_in_weight),
    .io_in_psum(PE_Array_6_2_io_in_psum),
    .io_in_flow(PE_Array_6_2_io_in_flow),
    .io_in_shift(PE_Array_6_2_io_in_shift),
    .io_out_activate(PE_Array_6_2_io_out_activate),
    .io_out_weight(PE_Array_6_2_io_out_weight),
    .io_out_psum(PE_Array_6_2_io_out_psum)
  );
  basic_PE PE_Array_6_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_3_clock),
    .reset(PE_Array_6_3_reset),
    .io_in_activate(PE_Array_6_3_io_in_activate),
    .io_in_weight(PE_Array_6_3_io_in_weight),
    .io_in_psum(PE_Array_6_3_io_in_psum),
    .io_in_flow(PE_Array_6_3_io_in_flow),
    .io_in_shift(PE_Array_6_3_io_in_shift),
    .io_out_activate(PE_Array_6_3_io_out_activate),
    .io_out_weight(PE_Array_6_3_io_out_weight),
    .io_out_psum(PE_Array_6_3_io_out_psum)
  );
  basic_PE PE_Array_6_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_4_clock),
    .reset(PE_Array_6_4_reset),
    .io_in_activate(PE_Array_6_4_io_in_activate),
    .io_in_weight(PE_Array_6_4_io_in_weight),
    .io_in_psum(PE_Array_6_4_io_in_psum),
    .io_in_flow(PE_Array_6_4_io_in_flow),
    .io_in_shift(PE_Array_6_4_io_in_shift),
    .io_out_activate(PE_Array_6_4_io_out_activate),
    .io_out_weight(PE_Array_6_4_io_out_weight),
    .io_out_psum(PE_Array_6_4_io_out_psum)
  );
  basic_PE PE_Array_6_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_5_clock),
    .reset(PE_Array_6_5_reset),
    .io_in_activate(PE_Array_6_5_io_in_activate),
    .io_in_weight(PE_Array_6_5_io_in_weight),
    .io_in_psum(PE_Array_6_5_io_in_psum),
    .io_in_flow(PE_Array_6_5_io_in_flow),
    .io_in_shift(PE_Array_6_5_io_in_shift),
    .io_out_activate(PE_Array_6_5_io_out_activate),
    .io_out_weight(PE_Array_6_5_io_out_weight),
    .io_out_psum(PE_Array_6_5_io_out_psum)
  );
  basic_PE PE_Array_6_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_6_clock),
    .reset(PE_Array_6_6_reset),
    .io_in_activate(PE_Array_6_6_io_in_activate),
    .io_in_weight(PE_Array_6_6_io_in_weight),
    .io_in_psum(PE_Array_6_6_io_in_psum),
    .io_in_flow(PE_Array_6_6_io_in_flow),
    .io_in_shift(PE_Array_6_6_io_in_shift),
    .io_out_activate(PE_Array_6_6_io_out_activate),
    .io_out_weight(PE_Array_6_6_io_out_weight),
    .io_out_psum(PE_Array_6_6_io_out_psum)
  );
  basic_PE PE_Array_6_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_6_7_clock),
    .reset(PE_Array_6_7_reset),
    .io_in_activate(PE_Array_6_7_io_in_activate),
    .io_in_weight(PE_Array_6_7_io_in_weight),
    .io_in_psum(PE_Array_6_7_io_in_psum),
    .io_in_flow(PE_Array_6_7_io_in_flow),
    .io_in_shift(PE_Array_6_7_io_in_shift),
    .io_out_activate(PE_Array_6_7_io_out_activate),
    .io_out_weight(PE_Array_6_7_io_out_weight),
    .io_out_psum(PE_Array_6_7_io_out_psum)
  );
  basic_PE PE_Array_7_0 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_0_clock),
    .reset(PE_Array_7_0_reset),
    .io_in_activate(PE_Array_7_0_io_in_activate),
    .io_in_weight(PE_Array_7_0_io_in_weight),
    .io_in_psum(PE_Array_7_0_io_in_psum),
    .io_in_flow(PE_Array_7_0_io_in_flow),
    .io_in_shift(PE_Array_7_0_io_in_shift),
    .io_out_activate(PE_Array_7_0_io_out_activate),
    .io_out_weight(PE_Array_7_0_io_out_weight),
    .io_out_psum(PE_Array_7_0_io_out_psum)
  );
  basic_PE PE_Array_7_1 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_1_clock),
    .reset(PE_Array_7_1_reset),
    .io_in_activate(PE_Array_7_1_io_in_activate),
    .io_in_weight(PE_Array_7_1_io_in_weight),
    .io_in_psum(PE_Array_7_1_io_in_psum),
    .io_in_flow(PE_Array_7_1_io_in_flow),
    .io_in_shift(PE_Array_7_1_io_in_shift),
    .io_out_activate(PE_Array_7_1_io_out_activate),
    .io_out_weight(PE_Array_7_1_io_out_weight),
    .io_out_psum(PE_Array_7_1_io_out_psum)
  );
  basic_PE PE_Array_7_2 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_2_clock),
    .reset(PE_Array_7_2_reset),
    .io_in_activate(PE_Array_7_2_io_in_activate),
    .io_in_weight(PE_Array_7_2_io_in_weight),
    .io_in_psum(PE_Array_7_2_io_in_psum),
    .io_in_flow(PE_Array_7_2_io_in_flow),
    .io_in_shift(PE_Array_7_2_io_in_shift),
    .io_out_activate(PE_Array_7_2_io_out_activate),
    .io_out_weight(PE_Array_7_2_io_out_weight),
    .io_out_psum(PE_Array_7_2_io_out_psum)
  );
  basic_PE PE_Array_7_3 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_3_clock),
    .reset(PE_Array_7_3_reset),
    .io_in_activate(PE_Array_7_3_io_in_activate),
    .io_in_weight(PE_Array_7_3_io_in_weight),
    .io_in_psum(PE_Array_7_3_io_in_psum),
    .io_in_flow(PE_Array_7_3_io_in_flow),
    .io_in_shift(PE_Array_7_3_io_in_shift),
    .io_out_activate(PE_Array_7_3_io_out_activate),
    .io_out_weight(PE_Array_7_3_io_out_weight),
    .io_out_psum(PE_Array_7_3_io_out_psum)
  );
  basic_PE PE_Array_7_4 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_4_clock),
    .reset(PE_Array_7_4_reset),
    .io_in_activate(PE_Array_7_4_io_in_activate),
    .io_in_weight(PE_Array_7_4_io_in_weight),
    .io_in_psum(PE_Array_7_4_io_in_psum),
    .io_in_flow(PE_Array_7_4_io_in_flow),
    .io_in_shift(PE_Array_7_4_io_in_shift),
    .io_out_activate(PE_Array_7_4_io_out_activate),
    .io_out_weight(PE_Array_7_4_io_out_weight),
    .io_out_psum(PE_Array_7_4_io_out_psum)
  );
  basic_PE PE_Array_7_5 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_5_clock),
    .reset(PE_Array_7_5_reset),
    .io_in_activate(PE_Array_7_5_io_in_activate),
    .io_in_weight(PE_Array_7_5_io_in_weight),
    .io_in_psum(PE_Array_7_5_io_in_psum),
    .io_in_flow(PE_Array_7_5_io_in_flow),
    .io_in_shift(PE_Array_7_5_io_in_shift),
    .io_out_activate(PE_Array_7_5_io_out_activate),
    .io_out_weight(PE_Array_7_5_io_out_weight),
    .io_out_psum(PE_Array_7_5_io_out_psum)
  );
  basic_PE PE_Array_7_6 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_6_clock),
    .reset(PE_Array_7_6_reset),
    .io_in_activate(PE_Array_7_6_io_in_activate),
    .io_in_weight(PE_Array_7_6_io_in_weight),
    .io_in_psum(PE_Array_7_6_io_in_psum),
    .io_in_flow(PE_Array_7_6_io_in_flow),
    .io_in_shift(PE_Array_7_6_io_in_shift),
    .io_out_activate(PE_Array_7_6_io_out_activate),
    .io_out_weight(PE_Array_7_6_io_out_weight),
    .io_out_psum(PE_Array_7_6_io_out_psum)
  );
  basic_PE PE_Array_7_7 ( // @[Systolic_Array.scala 19:62]
    .clock(PE_Array_7_7_clock),
    .reset(PE_Array_7_7_reset),
    .io_in_activate(PE_Array_7_7_io_in_activate),
    .io_in_weight(PE_Array_7_7_io_in_weight),
    .io_in_psum(PE_Array_7_7_io_in_psum),
    .io_in_flow(PE_Array_7_7_io_in_flow),
    .io_in_shift(PE_Array_7_7_io_in_shift),
    .io_out_activate(PE_Array_7_7_io_out_activate),
    .io_out_weight(PE_Array_7_7_io_out_weight),
    .io_out_psum(PE_Array_7_7_io_out_psum)
  );
  assign io_psum_0 = PE_Array_7_0_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_1 = PE_Array_7_1_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_2 = PE_Array_7_2_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_3 = PE_Array_7_3_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_4 = PE_Array_7_4_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_5 = PE_Array_7_5_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_6 = PE_Array_7_6_io_out_psum; // @[DataPath.scala 24:10]
  assign io_psum_7 = PE_Array_7_7_io_out_psum; // @[DataPath.scala 24:10]
  assign io_valid_0 = valid_reg[0]; // @[Systolic_Array.scala 73:33]
  assign io_valid_1 = valid_reg[1]; // @[Systolic_Array.scala 73:33]
  assign io_valid_2 = valid_reg[2]; // @[Systolic_Array.scala 73:33]
  assign io_valid_3 = valid_reg[3]; // @[Systolic_Array.scala 73:33]
  assign io_valid_4 = valid_reg[4]; // @[Systolic_Array.scala 73:33]
  assign io_valid_5 = valid_reg[5]; // @[Systolic_Array.scala 73:33]
  assign io_valid_6 = valid_reg[6]; // @[Systolic_Array.scala 73:33]
  assign io_valid_7 = valid_reg[7]; // @[Systolic_Array.scala 73:33]
  assign PE_Array_0_0_clock = clock;
  assign PE_Array_0_0_reset = reset;
  assign PE_Array_0_0_io_in_activate = io_activate_0; // @[DataPath.scala 11:26]
  assign PE_Array_0_0_io_in_weight = io_weight_0; // @[DataPath.scala 20:23]
  assign PE_Array_0_0_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_1_clock = clock;
  assign PE_Array_0_1_reset = reset;
  assign PE_Array_0_1_io_in_activate = PE_Array_0_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_1_io_in_weight = io_weight_1; // @[DataPath.scala 20:23]
  assign PE_Array_0_1_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_2_clock = clock;
  assign PE_Array_0_2_reset = reset;
  assign PE_Array_0_2_io_in_activate = PE_Array_0_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_2_io_in_weight = io_weight_2; // @[DataPath.scala 20:23]
  assign PE_Array_0_2_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_3_clock = clock;
  assign PE_Array_0_3_reset = reset;
  assign PE_Array_0_3_io_in_activate = PE_Array_0_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_3_io_in_weight = io_weight_3; // @[DataPath.scala 20:23]
  assign PE_Array_0_3_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_4_clock = clock;
  assign PE_Array_0_4_reset = reset;
  assign PE_Array_0_4_io_in_activate = PE_Array_0_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_4_io_in_weight = io_weight_4; // @[DataPath.scala 20:23]
  assign PE_Array_0_4_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_5_clock = clock;
  assign PE_Array_0_5_reset = reset;
  assign PE_Array_0_5_io_in_activate = PE_Array_0_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_5_io_in_weight = io_weight_5; // @[DataPath.scala 20:23]
  assign PE_Array_0_5_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_6_clock = clock;
  assign PE_Array_0_6_reset = reset;
  assign PE_Array_0_6_io_in_activate = PE_Array_0_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_6_io_in_weight = io_weight_6; // @[DataPath.scala 20:23]
  assign PE_Array_0_6_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_0_7_clock = clock;
  assign PE_Array_0_7_reset = reset;
  assign PE_Array_0_7_io_in_activate = PE_Array_0_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_0_7_io_in_weight = io_weight_7; // @[DataPath.scala 20:23]
  assign PE_Array_0_7_io_in_psum = 16'h0; // @[DataPath.scala 21:21]
  assign PE_Array_0_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_0_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_0_clock = clock;
  assign PE_Array_1_0_reset = reset;
  assign PE_Array_1_0_io_in_activate = io_activate_1; // @[DataPath.scala 11:26]
  assign PE_Array_1_0_io_in_weight = PE_Array_0_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_0_io_in_psum = PE_Array_0_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_1_clock = clock;
  assign PE_Array_1_1_reset = reset;
  assign PE_Array_1_1_io_in_activate = PE_Array_1_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_1_io_in_weight = PE_Array_0_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_1_io_in_psum = PE_Array_0_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_2_clock = clock;
  assign PE_Array_1_2_reset = reset;
  assign PE_Array_1_2_io_in_activate = PE_Array_1_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_2_io_in_weight = PE_Array_0_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_2_io_in_psum = PE_Array_0_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_3_clock = clock;
  assign PE_Array_1_3_reset = reset;
  assign PE_Array_1_3_io_in_activate = PE_Array_1_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_3_io_in_weight = PE_Array_0_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_3_io_in_psum = PE_Array_0_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_4_clock = clock;
  assign PE_Array_1_4_reset = reset;
  assign PE_Array_1_4_io_in_activate = PE_Array_1_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_4_io_in_weight = PE_Array_0_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_4_io_in_psum = PE_Array_0_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_5_clock = clock;
  assign PE_Array_1_5_reset = reset;
  assign PE_Array_1_5_io_in_activate = PE_Array_1_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_5_io_in_weight = PE_Array_0_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_5_io_in_psum = PE_Array_0_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_6_clock = clock;
  assign PE_Array_1_6_reset = reset;
  assign PE_Array_1_6_io_in_activate = PE_Array_1_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_6_io_in_weight = PE_Array_0_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_6_io_in_psum = PE_Array_0_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_1_7_clock = clock;
  assign PE_Array_1_7_reset = reset;
  assign PE_Array_1_7_io_in_activate = PE_Array_1_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_1_7_io_in_weight = PE_Array_0_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_1_7_io_in_psum = PE_Array_0_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_1_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_1_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_0_clock = clock;
  assign PE_Array_2_0_reset = reset;
  assign PE_Array_2_0_io_in_activate = io_activate_2; // @[DataPath.scala 11:26]
  assign PE_Array_2_0_io_in_weight = PE_Array_1_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_0_io_in_psum = PE_Array_1_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_1_clock = clock;
  assign PE_Array_2_1_reset = reset;
  assign PE_Array_2_1_io_in_activate = PE_Array_2_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_1_io_in_weight = PE_Array_1_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_1_io_in_psum = PE_Array_1_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_2_clock = clock;
  assign PE_Array_2_2_reset = reset;
  assign PE_Array_2_2_io_in_activate = PE_Array_2_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_2_io_in_weight = PE_Array_1_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_2_io_in_psum = PE_Array_1_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_3_clock = clock;
  assign PE_Array_2_3_reset = reset;
  assign PE_Array_2_3_io_in_activate = PE_Array_2_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_3_io_in_weight = PE_Array_1_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_3_io_in_psum = PE_Array_1_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_4_clock = clock;
  assign PE_Array_2_4_reset = reset;
  assign PE_Array_2_4_io_in_activate = PE_Array_2_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_4_io_in_weight = PE_Array_1_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_4_io_in_psum = PE_Array_1_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_5_clock = clock;
  assign PE_Array_2_5_reset = reset;
  assign PE_Array_2_5_io_in_activate = PE_Array_2_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_5_io_in_weight = PE_Array_1_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_5_io_in_psum = PE_Array_1_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_6_clock = clock;
  assign PE_Array_2_6_reset = reset;
  assign PE_Array_2_6_io_in_activate = PE_Array_2_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_6_io_in_weight = PE_Array_1_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_6_io_in_psum = PE_Array_1_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_2_7_clock = clock;
  assign PE_Array_2_7_reset = reset;
  assign PE_Array_2_7_io_in_activate = PE_Array_2_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_2_7_io_in_weight = PE_Array_1_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_2_7_io_in_psum = PE_Array_1_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_2_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_2_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_0_clock = clock;
  assign PE_Array_3_0_reset = reset;
  assign PE_Array_3_0_io_in_activate = io_activate_3; // @[DataPath.scala 11:26]
  assign PE_Array_3_0_io_in_weight = PE_Array_2_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_0_io_in_psum = PE_Array_2_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_1_clock = clock;
  assign PE_Array_3_1_reset = reset;
  assign PE_Array_3_1_io_in_activate = PE_Array_3_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_1_io_in_weight = PE_Array_2_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_1_io_in_psum = PE_Array_2_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_2_clock = clock;
  assign PE_Array_3_2_reset = reset;
  assign PE_Array_3_2_io_in_activate = PE_Array_3_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_2_io_in_weight = PE_Array_2_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_2_io_in_psum = PE_Array_2_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_3_clock = clock;
  assign PE_Array_3_3_reset = reset;
  assign PE_Array_3_3_io_in_activate = PE_Array_3_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_3_io_in_weight = PE_Array_2_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_3_io_in_psum = PE_Array_2_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_4_clock = clock;
  assign PE_Array_3_4_reset = reset;
  assign PE_Array_3_4_io_in_activate = PE_Array_3_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_4_io_in_weight = PE_Array_2_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_4_io_in_psum = PE_Array_2_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_5_clock = clock;
  assign PE_Array_3_5_reset = reset;
  assign PE_Array_3_5_io_in_activate = PE_Array_3_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_5_io_in_weight = PE_Array_2_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_5_io_in_psum = PE_Array_2_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_6_clock = clock;
  assign PE_Array_3_6_reset = reset;
  assign PE_Array_3_6_io_in_activate = PE_Array_3_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_6_io_in_weight = PE_Array_2_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_6_io_in_psum = PE_Array_2_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_3_7_clock = clock;
  assign PE_Array_3_7_reset = reset;
  assign PE_Array_3_7_io_in_activate = PE_Array_3_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_3_7_io_in_weight = PE_Array_2_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_3_7_io_in_psum = PE_Array_2_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_3_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_3_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_0_clock = clock;
  assign PE_Array_4_0_reset = reset;
  assign PE_Array_4_0_io_in_activate = io_activate_4; // @[DataPath.scala 11:26]
  assign PE_Array_4_0_io_in_weight = PE_Array_3_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_0_io_in_psum = PE_Array_3_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_1_clock = clock;
  assign PE_Array_4_1_reset = reset;
  assign PE_Array_4_1_io_in_activate = PE_Array_4_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_1_io_in_weight = PE_Array_3_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_1_io_in_psum = PE_Array_3_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_2_clock = clock;
  assign PE_Array_4_2_reset = reset;
  assign PE_Array_4_2_io_in_activate = PE_Array_4_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_2_io_in_weight = PE_Array_3_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_2_io_in_psum = PE_Array_3_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_3_clock = clock;
  assign PE_Array_4_3_reset = reset;
  assign PE_Array_4_3_io_in_activate = PE_Array_4_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_3_io_in_weight = PE_Array_3_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_3_io_in_psum = PE_Array_3_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_4_clock = clock;
  assign PE_Array_4_4_reset = reset;
  assign PE_Array_4_4_io_in_activate = PE_Array_4_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_4_io_in_weight = PE_Array_3_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_4_io_in_psum = PE_Array_3_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_5_clock = clock;
  assign PE_Array_4_5_reset = reset;
  assign PE_Array_4_5_io_in_activate = PE_Array_4_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_5_io_in_weight = PE_Array_3_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_5_io_in_psum = PE_Array_3_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_6_clock = clock;
  assign PE_Array_4_6_reset = reset;
  assign PE_Array_4_6_io_in_activate = PE_Array_4_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_6_io_in_weight = PE_Array_3_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_6_io_in_psum = PE_Array_3_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_4_7_clock = clock;
  assign PE_Array_4_7_reset = reset;
  assign PE_Array_4_7_io_in_activate = PE_Array_4_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_4_7_io_in_weight = PE_Array_3_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_4_7_io_in_psum = PE_Array_3_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_4_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_4_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_0_clock = clock;
  assign PE_Array_5_0_reset = reset;
  assign PE_Array_5_0_io_in_activate = io_activate_5; // @[DataPath.scala 11:26]
  assign PE_Array_5_0_io_in_weight = PE_Array_4_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_0_io_in_psum = PE_Array_4_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_1_clock = clock;
  assign PE_Array_5_1_reset = reset;
  assign PE_Array_5_1_io_in_activate = PE_Array_5_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_1_io_in_weight = PE_Array_4_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_1_io_in_psum = PE_Array_4_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_2_clock = clock;
  assign PE_Array_5_2_reset = reset;
  assign PE_Array_5_2_io_in_activate = PE_Array_5_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_2_io_in_weight = PE_Array_4_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_2_io_in_psum = PE_Array_4_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_3_clock = clock;
  assign PE_Array_5_3_reset = reset;
  assign PE_Array_5_3_io_in_activate = PE_Array_5_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_3_io_in_weight = PE_Array_4_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_3_io_in_psum = PE_Array_4_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_4_clock = clock;
  assign PE_Array_5_4_reset = reset;
  assign PE_Array_5_4_io_in_activate = PE_Array_5_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_4_io_in_weight = PE_Array_4_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_4_io_in_psum = PE_Array_4_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_5_clock = clock;
  assign PE_Array_5_5_reset = reset;
  assign PE_Array_5_5_io_in_activate = PE_Array_5_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_5_io_in_weight = PE_Array_4_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_5_io_in_psum = PE_Array_4_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_6_clock = clock;
  assign PE_Array_5_6_reset = reset;
  assign PE_Array_5_6_io_in_activate = PE_Array_5_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_6_io_in_weight = PE_Array_4_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_6_io_in_psum = PE_Array_4_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_5_7_clock = clock;
  assign PE_Array_5_7_reset = reset;
  assign PE_Array_5_7_io_in_activate = PE_Array_5_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_5_7_io_in_weight = PE_Array_4_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_5_7_io_in_psum = PE_Array_4_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_5_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_5_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_0_clock = clock;
  assign PE_Array_6_0_reset = reset;
  assign PE_Array_6_0_io_in_activate = io_activate_6; // @[DataPath.scala 11:26]
  assign PE_Array_6_0_io_in_weight = PE_Array_5_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_0_io_in_psum = PE_Array_5_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_1_clock = clock;
  assign PE_Array_6_1_reset = reset;
  assign PE_Array_6_1_io_in_activate = PE_Array_6_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_1_io_in_weight = PE_Array_5_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_1_io_in_psum = PE_Array_5_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_2_clock = clock;
  assign PE_Array_6_2_reset = reset;
  assign PE_Array_6_2_io_in_activate = PE_Array_6_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_2_io_in_weight = PE_Array_5_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_2_io_in_psum = PE_Array_5_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_3_clock = clock;
  assign PE_Array_6_3_reset = reset;
  assign PE_Array_6_3_io_in_activate = PE_Array_6_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_3_io_in_weight = PE_Array_5_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_3_io_in_psum = PE_Array_5_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_4_clock = clock;
  assign PE_Array_6_4_reset = reset;
  assign PE_Array_6_4_io_in_activate = PE_Array_6_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_4_io_in_weight = PE_Array_5_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_4_io_in_psum = PE_Array_5_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_5_clock = clock;
  assign PE_Array_6_5_reset = reset;
  assign PE_Array_6_5_io_in_activate = PE_Array_6_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_5_io_in_weight = PE_Array_5_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_5_io_in_psum = PE_Array_5_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_6_clock = clock;
  assign PE_Array_6_6_reset = reset;
  assign PE_Array_6_6_io_in_activate = PE_Array_6_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_6_io_in_weight = PE_Array_5_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_6_io_in_psum = PE_Array_5_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_6_7_clock = clock;
  assign PE_Array_6_7_reset = reset;
  assign PE_Array_6_7_io_in_activate = PE_Array_6_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_6_7_io_in_weight = PE_Array_5_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_6_7_io_in_psum = PE_Array_5_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_6_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_6_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_0_clock = clock;
  assign PE_Array_7_0_reset = reset;
  assign PE_Array_7_0_io_in_activate = io_activate_7; // @[DataPath.scala 11:26]
  assign PE_Array_7_0_io_in_weight = PE_Array_6_0_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_0_io_in_psum = PE_Array_6_0_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_0_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_0_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_1_clock = clock;
  assign PE_Array_7_1_reset = reset;
  assign PE_Array_7_1_io_in_activate = PE_Array_7_0_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_1_io_in_weight = PE_Array_6_1_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_1_io_in_psum = PE_Array_6_1_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_1_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_1_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_2_clock = clock;
  assign PE_Array_7_2_reset = reset;
  assign PE_Array_7_2_io_in_activate = PE_Array_7_1_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_2_io_in_weight = PE_Array_6_2_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_2_io_in_psum = PE_Array_6_2_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_2_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_2_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_3_clock = clock;
  assign PE_Array_7_3_reset = reset;
  assign PE_Array_7_3_io_in_activate = PE_Array_7_2_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_3_io_in_weight = PE_Array_6_3_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_3_io_in_psum = PE_Array_6_3_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_3_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_3_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_4_clock = clock;
  assign PE_Array_7_4_reset = reset;
  assign PE_Array_7_4_io_in_activate = PE_Array_7_3_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_4_io_in_weight = PE_Array_6_4_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_4_io_in_psum = PE_Array_6_4_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_4_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_4_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_5_clock = clock;
  assign PE_Array_7_5_reset = reset;
  assign PE_Array_7_5_io_in_activate = PE_Array_7_4_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_5_io_in_weight = PE_Array_6_5_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_5_io_in_psum = PE_Array_6_5_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_5_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_5_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_6_clock = clock;
  assign PE_Array_7_6_reset = reset;
  assign PE_Array_7_6_io_in_activate = PE_Array_7_5_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_6_io_in_weight = PE_Array_6_6_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_6_io_in_psum = PE_Array_6_6_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_6_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_6_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  assign PE_Array_7_7_clock = clock;
  assign PE_Array_7_7_reset = reset;
  assign PE_Array_7_7_io_in_activate = PE_Array_7_6_io_out_activate; // @[DataPath.scala 7:26]
  assign PE_Array_7_7_io_in_weight = PE_Array_6_7_io_out_weight; // @[DataPath.scala 15:23]
  assign PE_Array_7_7_io_in_psum = PE_Array_6_7_io_out_psum; // @[DataPath.scala 16:21]
  assign PE_Array_7_7_io_in_flow = io_flow; // @[Systolic_Array.scala 22:54]
  assign PE_Array_7_7_io_in_shift = io_shift; // @[Systolic_Array.scala 23:55]
  always @(posedge clock) begin
    if (reset) begin // @[Systolic_Array.scala 52:29]
      flow_counter <= 5'h0; // @[Systolic_Array.scala 52:29]
    end else if (io_flow & flow_counter < 5'h16) begin // @[Systolic_Array.scala 56:58]
      flow_counter <= _flow_counter_T_1; // @[Systolic_Array.scala 57:18]
    end else if (flow_counter == 5'h16) begin // @[Systolic_Array.scala 58:53]
      flow_counter <= 5'h0; // @[Systolic_Array.scala 59:18]
    end
    if (reset) begin // @[Systolic_Array.scala 53:26]
      valid_reg <= 8'h0; // @[Systolic_Array.scala 53:26]
    end else if (io_flow & 5'h7 <= flow_counter & flow_counter < 5'hf) begin // @[Systolic_Array.scala 65:96]
      valid_reg <= _valid_reg_T_1; // @[Systolic_Array.scala 66:15]
    end else if (io_flow & flow_counter >= 5'hf) begin // @[Systolic_Array.scala 67:65]
      valid_reg <= _valid_reg_T_3; // @[Systolic_Array.scala 68:15]
    end else begin
      valid_reg <= 8'h0; // @[Systolic_Array.scala 70:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flow_counter = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Accumulator_Array(
  input         clock,
  input         reset,
  input  [15:0] io_in_psum_0,
  input  [15:0] io_in_psum_1,
  input  [15:0] io_in_psum_2,
  input  [15:0] io_in_psum_3,
  input  [15:0] io_in_psum_4,
  input  [15:0] io_in_psum_5,
  input  [15:0] io_in_psum_6,
  input  [15:0] io_in_psum_7,
  input         io_in_valid_0,
  input         io_in_valid_1,
  input         io_in_valid_2,
  input         io_in_valid_3,
  input         io_in_valid_4,
  input         io_in_valid_5,
  input         io_in_valid_6,
  input         io_in_valid_7,
  input         io_in_acc,
  input         io_in_compute_done,
  output        io_isdone,
  output [31:0] io_out_sum_0,
  output [31:0] io_out_sum_1,
  output [31:0] io_out_sum_2,
  output [31:0] io_out_sum_3,
  output [31:0] io_out_sum_4,
  output [31:0] io_out_sum_5,
  output [31:0] io_out_sum_6,
  output [31:0] io_out_sum_7,
  output [31:0] io_out_sum_8,
  output [31:0] io_out_sum_9,
  output [31:0] io_out_sum_10,
  output [31:0] io_out_sum_11,
  output [31:0] io_out_sum_12,
  output [31:0] io_out_sum_13,
  output [31:0] io_out_sum_14,
  output [31:0] io_out_sum_15,
  output [31:0] io_out_sum_16,
  output [31:0] io_out_sum_17,
  output [31:0] io_out_sum_18,
  output [31:0] io_out_sum_19,
  output [31:0] io_out_sum_20,
  output [31:0] io_out_sum_21,
  output [31:0] io_out_sum_22,
  output [31:0] io_out_sum_23,
  output [31:0] io_out_sum_24,
  output [31:0] io_out_sum_25,
  output [31:0] io_out_sum_26,
  output [31:0] io_out_sum_27,
  output [31:0] io_out_sum_28,
  output [31:0] io_out_sum_29,
  output [31:0] io_out_sum_30,
  output [31:0] io_out_sum_31,
  output [31:0] io_out_sum_32,
  output [31:0] io_out_sum_33,
  output [31:0] io_out_sum_34,
  output [31:0] io_out_sum_35,
  output [31:0] io_out_sum_36,
  output [31:0] io_out_sum_37,
  output [31:0] io_out_sum_38,
  output [31:0] io_out_sum_39,
  output [31:0] io_out_sum_40,
  output [31:0] io_out_sum_41,
  output [31:0] io_out_sum_42,
  output [31:0] io_out_sum_43,
  output [31:0] io_out_sum_44,
  output [31:0] io_out_sum_45,
  output [31:0] io_out_sum_46,
  output [31:0] io_out_sum_47,
  output [31:0] io_out_sum_48,
  output [31:0] io_out_sum_49,
  output [31:0] io_out_sum_50,
  output [31:0] io_out_sum_51,
  output [31:0] io_out_sum_52,
  output [31:0] io_out_sum_53,
  output [31:0] io_out_sum_54,
  output [31:0] io_out_sum_55,
  output [31:0] io_out_sum_56,
  output [31:0] io_out_sum_57,
  output [31:0] io_out_sum_58,
  output [31:0] io_out_sum_59,
  output [31:0] io_out_sum_60,
  output [31:0] io_out_sum_61,
  output [31:0] io_out_sum_62,
  output [31:0] io_out_sum_63,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] Acc_Buffer_0_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_0_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_1_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_2_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_3_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_4_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_5_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_6_7; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_0; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_1; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_2; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_3; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_4; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_5; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_6; // @[Accumulator_Array.scala 20:27]
  reg [15:0] Acc_Buffer_7_7; // @[Accumulator_Array.scala 20:27]
  reg [31:0] Acc_Result_0_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_0_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_1_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_2_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_3_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_4_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_5_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_6_7; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_0; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_1; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_2; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_3; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_4; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_5; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_6; // @[Accumulator_Array.scala 21:27]
  reg [31:0] Acc_Result_7_7; // @[Accumulator_Array.scala 21:27]
  reg [3:0] valid_counter_0; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_1; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_2; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_3; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_4; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_5; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_6; // @[Accumulator_Array.scala 22:30]
  reg [3:0] valid_counter_7; // @[Accumulator_Array.scala 22:30]
  wire [15:0] _GEN_17 = 3'h1 == valid_counter_0[2:0] ? Acc_Buffer_1_0 : Acc_Buffer_0_0; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_18 = 3'h2 == valid_counter_0[2:0] ? Acc_Buffer_2_0 : _GEN_17; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_19 = 3'h3 == valid_counter_0[2:0] ? Acc_Buffer_3_0 : _GEN_18; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_20 = 3'h4 == valid_counter_0[2:0] ? Acc_Buffer_4_0 : _GEN_19; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_21 = 3'h5 == valid_counter_0[2:0] ? Acc_Buffer_5_0 : _GEN_20; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_22 = 3'h6 == valid_counter_0[2:0] ? Acc_Buffer_6_0 : _GEN_21; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_49 = 3'h1 == valid_counter_1[2:0] ? Acc_Buffer_1_1 : Acc_Buffer_0_1; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_50 = 3'h2 == valid_counter_1[2:0] ? Acc_Buffer_2_1 : _GEN_49; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_51 = 3'h3 == valid_counter_1[2:0] ? Acc_Buffer_3_1 : _GEN_50; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_52 = 3'h4 == valid_counter_1[2:0] ? Acc_Buffer_4_1 : _GEN_51; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_53 = 3'h5 == valid_counter_1[2:0] ? Acc_Buffer_5_1 : _GEN_52; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_54 = 3'h6 == valid_counter_1[2:0] ? Acc_Buffer_6_1 : _GEN_53; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_81 = 3'h1 == valid_counter_2[2:0] ? Acc_Buffer_1_2 : Acc_Buffer_0_2; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_82 = 3'h2 == valid_counter_2[2:0] ? Acc_Buffer_2_2 : _GEN_81; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_83 = 3'h3 == valid_counter_2[2:0] ? Acc_Buffer_3_2 : _GEN_82; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_84 = 3'h4 == valid_counter_2[2:0] ? Acc_Buffer_4_2 : _GEN_83; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_85 = 3'h5 == valid_counter_2[2:0] ? Acc_Buffer_5_2 : _GEN_84; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_86 = 3'h6 == valid_counter_2[2:0] ? Acc_Buffer_6_2 : _GEN_85; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_113 = 3'h1 == valid_counter_3[2:0] ? Acc_Buffer_1_3 : Acc_Buffer_0_3; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_114 = 3'h2 == valid_counter_3[2:0] ? Acc_Buffer_2_3 : _GEN_113; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_115 = 3'h3 == valid_counter_3[2:0] ? Acc_Buffer_3_3 : _GEN_114; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_116 = 3'h4 == valid_counter_3[2:0] ? Acc_Buffer_4_3 : _GEN_115; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_117 = 3'h5 == valid_counter_3[2:0] ? Acc_Buffer_5_3 : _GEN_116; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_118 = 3'h6 == valid_counter_3[2:0] ? Acc_Buffer_6_3 : _GEN_117; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_145 = 3'h1 == valid_counter_4[2:0] ? Acc_Buffer_1_4 : Acc_Buffer_0_4; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_146 = 3'h2 == valid_counter_4[2:0] ? Acc_Buffer_2_4 : _GEN_145; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_147 = 3'h3 == valid_counter_4[2:0] ? Acc_Buffer_3_4 : _GEN_146; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_148 = 3'h4 == valid_counter_4[2:0] ? Acc_Buffer_4_4 : _GEN_147; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_149 = 3'h5 == valid_counter_4[2:0] ? Acc_Buffer_5_4 : _GEN_148; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_150 = 3'h6 == valid_counter_4[2:0] ? Acc_Buffer_6_4 : _GEN_149; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_177 = 3'h1 == valid_counter_5[2:0] ? Acc_Buffer_1_5 : Acc_Buffer_0_5; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_178 = 3'h2 == valid_counter_5[2:0] ? Acc_Buffer_2_5 : _GEN_177; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_179 = 3'h3 == valid_counter_5[2:0] ? Acc_Buffer_3_5 : _GEN_178; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_180 = 3'h4 == valid_counter_5[2:0] ? Acc_Buffer_4_5 : _GEN_179; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_181 = 3'h5 == valid_counter_5[2:0] ? Acc_Buffer_5_5 : _GEN_180; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_182 = 3'h6 == valid_counter_5[2:0] ? Acc_Buffer_6_5 : _GEN_181; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_209 = 3'h1 == valid_counter_6[2:0] ? Acc_Buffer_1_6 : Acc_Buffer_0_6; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_210 = 3'h2 == valid_counter_6[2:0] ? Acc_Buffer_2_6 : _GEN_209; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_211 = 3'h3 == valid_counter_6[2:0] ? Acc_Buffer_3_6 : _GEN_210; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_212 = 3'h4 == valid_counter_6[2:0] ? Acc_Buffer_4_6 : _GEN_211; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_213 = 3'h5 == valid_counter_6[2:0] ? Acc_Buffer_5_6 : _GEN_212; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_214 = 3'h6 == valid_counter_6[2:0] ? Acc_Buffer_6_6 : _GEN_213; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_241 = 3'h1 == valid_counter_7[2:0] ? Acc_Buffer_1_7 : Acc_Buffer_0_7; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_242 = 3'h2 == valid_counter_7[2:0] ? Acc_Buffer_2_7 : _GEN_241; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_243 = 3'h3 == valid_counter_7[2:0] ? Acc_Buffer_3_7 : _GEN_242; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_244 = 3'h4 == valid_counter_7[2:0] ? Acc_Buffer_4_7 : _GEN_243; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_245 = 3'h5 == valid_counter_7[2:0] ? Acc_Buffer_5_7 : _GEN_244; // @[Accumulator_Array.scala 28:{39,39}]
  wire [15:0] _GEN_246 = 3'h6 == valid_counter_7[2:0] ? Acc_Buffer_6_7 : _GEN_245; // @[Accumulator_Array.scala 28:{39,39}]
  wire [3:0] _valid_counter_0_T_1 = valid_counter_0 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_1_T_1 = valid_counter_1 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_2_T_1 = valid_counter_2 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_3_T_1 = valid_counter_3 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_4_T_1 = valid_counter_4 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_5_T_1 = valid_counter_5 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_6_T_1 = valid_counter_6 + 4'h1; // @[Accumulator_Array.scala 35:44]
  wire [3:0] _valid_counter_7_T_1 = valid_counter_7 + 4'h1; // @[Accumulator_Array.scala 35:44]
  reg [3:0] acc_counter; // @[Accumulator_Array.scala 43:28]
  wire [3:0] _acc_counter_T_1 = acc_counter + 4'h1; // @[Accumulator_Array.scala 46:32]
  wire  _T_43 = acc_counter != 4'h0; // @[Accumulator_Array.scala 49:26]
  wire [3:0] _T_46 = acc_counter - 4'h1; // @[Accumulator_Array.scala 57:30]
  wire [31:0] _GEN_276 = 3'h1 == _T_46[2:0] ? Acc_Result_1_0 : Acc_Result_0_0; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_277 = 3'h2 == _T_46[2:0] ? Acc_Result_2_0 : _GEN_276; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_278 = 3'h3 == _T_46[2:0] ? Acc_Result_3_0 : _GEN_277; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_279 = 3'h4 == _T_46[2:0] ? Acc_Result_4_0 : _GEN_278; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_280 = 3'h5 == _T_46[2:0] ? Acc_Result_5_0 : _GEN_279; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_281 = 3'h6 == _T_46[2:0] ? Acc_Result_6_0 : _GEN_280; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_282 = 3'h7 == _T_46[2:0] ? Acc_Result_7_0 : _GEN_281; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_284 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_0 : Acc_Buffer_0_0; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_285 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_0 : _GEN_284; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_286 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_0 : _GEN_285; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_287 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_0 : _GEN_286; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_288 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_0 : _GEN_287; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_289 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_0 : _GEN_288; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_290 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_0 : _GEN_289; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_597 = {{16'd0}, _GEN_290}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_0_T_7 = _GEN_282 + _GEN_597; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_300 = 3'h1 == _T_46[2:0] ? Acc_Result_1_1 : Acc_Result_0_1; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_301 = 3'h2 == _T_46[2:0] ? Acc_Result_2_1 : _GEN_300; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_302 = 3'h3 == _T_46[2:0] ? Acc_Result_3_1 : _GEN_301; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_303 = 3'h4 == _T_46[2:0] ? Acc_Result_4_1 : _GEN_302; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_304 = 3'h5 == _T_46[2:0] ? Acc_Result_5_1 : _GEN_303; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_305 = 3'h6 == _T_46[2:0] ? Acc_Result_6_1 : _GEN_304; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_306 = 3'h7 == _T_46[2:0] ? Acc_Result_7_1 : _GEN_305; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_308 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_1 : Acc_Buffer_0_1; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_309 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_1 : _GEN_308; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_310 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_1 : _GEN_309; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_311 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_1 : _GEN_310; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_312 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_1 : _GEN_311; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_313 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_1 : _GEN_312; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_314 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_1 : _GEN_313; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_598 = {{16'd0}, _GEN_314}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_1_T_7 = _GEN_306 + _GEN_598; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_324 = 3'h1 == _T_46[2:0] ? Acc_Result_1_2 : Acc_Result_0_2; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_325 = 3'h2 == _T_46[2:0] ? Acc_Result_2_2 : _GEN_324; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_326 = 3'h3 == _T_46[2:0] ? Acc_Result_3_2 : _GEN_325; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_327 = 3'h4 == _T_46[2:0] ? Acc_Result_4_2 : _GEN_326; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_328 = 3'h5 == _T_46[2:0] ? Acc_Result_5_2 : _GEN_327; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_329 = 3'h6 == _T_46[2:0] ? Acc_Result_6_2 : _GEN_328; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_330 = 3'h7 == _T_46[2:0] ? Acc_Result_7_2 : _GEN_329; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_332 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_2 : Acc_Buffer_0_2; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_333 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_2 : _GEN_332; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_334 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_2 : _GEN_333; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_335 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_2 : _GEN_334; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_336 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_2 : _GEN_335; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_337 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_2 : _GEN_336; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_338 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_2 : _GEN_337; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_599 = {{16'd0}, _GEN_338}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_2_T_7 = _GEN_330 + _GEN_599; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_348 = 3'h1 == _T_46[2:0] ? Acc_Result_1_3 : Acc_Result_0_3; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_349 = 3'h2 == _T_46[2:0] ? Acc_Result_2_3 : _GEN_348; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_350 = 3'h3 == _T_46[2:0] ? Acc_Result_3_3 : _GEN_349; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_351 = 3'h4 == _T_46[2:0] ? Acc_Result_4_3 : _GEN_350; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_352 = 3'h5 == _T_46[2:0] ? Acc_Result_5_3 : _GEN_351; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_353 = 3'h6 == _T_46[2:0] ? Acc_Result_6_3 : _GEN_352; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_354 = 3'h7 == _T_46[2:0] ? Acc_Result_7_3 : _GEN_353; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_356 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_3 : Acc_Buffer_0_3; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_357 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_3 : _GEN_356; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_358 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_3 : _GEN_357; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_359 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_3 : _GEN_358; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_360 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_3 : _GEN_359; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_361 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_3 : _GEN_360; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_362 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_3 : _GEN_361; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_600 = {{16'd0}, _GEN_362}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_3_T_7 = _GEN_354 + _GEN_600; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_372 = 3'h1 == _T_46[2:0] ? Acc_Result_1_4 : Acc_Result_0_4; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_373 = 3'h2 == _T_46[2:0] ? Acc_Result_2_4 : _GEN_372; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_374 = 3'h3 == _T_46[2:0] ? Acc_Result_3_4 : _GEN_373; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_375 = 3'h4 == _T_46[2:0] ? Acc_Result_4_4 : _GEN_374; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_376 = 3'h5 == _T_46[2:0] ? Acc_Result_5_4 : _GEN_375; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_377 = 3'h6 == _T_46[2:0] ? Acc_Result_6_4 : _GEN_376; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_378 = 3'h7 == _T_46[2:0] ? Acc_Result_7_4 : _GEN_377; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_380 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_4 : Acc_Buffer_0_4; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_381 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_4 : _GEN_380; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_382 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_4 : _GEN_381; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_383 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_4 : _GEN_382; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_384 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_4 : _GEN_383; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_385 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_4 : _GEN_384; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_386 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_4 : _GEN_385; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_601 = {{16'd0}, _GEN_386}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_4_T_7 = _GEN_378 + _GEN_601; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_396 = 3'h1 == _T_46[2:0] ? Acc_Result_1_5 : Acc_Result_0_5; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_397 = 3'h2 == _T_46[2:0] ? Acc_Result_2_5 : _GEN_396; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_398 = 3'h3 == _T_46[2:0] ? Acc_Result_3_5 : _GEN_397; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_399 = 3'h4 == _T_46[2:0] ? Acc_Result_4_5 : _GEN_398; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_400 = 3'h5 == _T_46[2:0] ? Acc_Result_5_5 : _GEN_399; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_401 = 3'h6 == _T_46[2:0] ? Acc_Result_6_5 : _GEN_400; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_402 = 3'h7 == _T_46[2:0] ? Acc_Result_7_5 : _GEN_401; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_404 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_5 : Acc_Buffer_0_5; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_405 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_5 : _GEN_404; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_406 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_5 : _GEN_405; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_407 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_5 : _GEN_406; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_408 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_5 : _GEN_407; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_409 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_5 : _GEN_408; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_410 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_5 : _GEN_409; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_602 = {{16'd0}, _GEN_410}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_5_T_7 = _GEN_402 + _GEN_602; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_420 = 3'h1 == _T_46[2:0] ? Acc_Result_1_6 : Acc_Result_0_6; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_421 = 3'h2 == _T_46[2:0] ? Acc_Result_2_6 : _GEN_420; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_422 = 3'h3 == _T_46[2:0] ? Acc_Result_3_6 : _GEN_421; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_423 = 3'h4 == _T_46[2:0] ? Acc_Result_4_6 : _GEN_422; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_424 = 3'h5 == _T_46[2:0] ? Acc_Result_5_6 : _GEN_423; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_425 = 3'h6 == _T_46[2:0] ? Acc_Result_6_6 : _GEN_424; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_426 = 3'h7 == _T_46[2:0] ? Acc_Result_7_6 : _GEN_425; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_428 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_6 : Acc_Buffer_0_6; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_429 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_6 : _GEN_428; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_430 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_6 : _GEN_429; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_431 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_6 : _GEN_430; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_432 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_6 : _GEN_431; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_433 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_6 : _GEN_432; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_434 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_6 : _GEN_433; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_603 = {{16'd0}, _GEN_434}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_6_T_7 = _GEN_426 + _GEN_603; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _GEN_444 = 3'h1 == _T_46[2:0] ? Acc_Result_1_7 : Acc_Result_0_7; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_445 = 3'h2 == _T_46[2:0] ? Acc_Result_2_7 : _GEN_444; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_446 = 3'h3 == _T_46[2:0] ? Acc_Result_3_7 : _GEN_445; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_447 = 3'h4 == _T_46[2:0] ? Acc_Result_4_7 : _GEN_446; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_448 = 3'h5 == _T_46[2:0] ? Acc_Result_5_7 : _GEN_447; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_449 = 3'h6 == _T_46[2:0] ? Acc_Result_6_7 : _GEN_448; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_450 = 3'h7 == _T_46[2:0] ? Acc_Result_7_7 : _GEN_449; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_452 = 3'h1 == _T_46[2:0] ? Acc_Buffer_1_7 : Acc_Buffer_0_7; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_453 = 3'h2 == _T_46[2:0] ? Acc_Buffer_2_7 : _GEN_452; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_454 = 3'h3 == _T_46[2:0] ? Acc_Buffer_3_7 : _GEN_453; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_455 = 3'h4 == _T_46[2:0] ? Acc_Buffer_4_7 : _GEN_454; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_456 = 3'h5 == _T_46[2:0] ? Acc_Buffer_5_7 : _GEN_455; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_457 = 3'h6 == _T_46[2:0] ? Acc_Buffer_6_7 : _GEN_456; // @[Accumulator_Array.scala 57:{76,76}]
  wire [15:0] _GEN_458 = 3'h7 == _T_46[2:0] ? Acc_Buffer_7_7 : _GEN_457; // @[Accumulator_Array.scala 57:{76,76}]
  wire [31:0] _GEN_604 = {{16'd0}, _GEN_458}; // @[Accumulator_Array.scala 57:76]
  wire [31:0] _Acc_Result_7_T_7 = _GEN_450 + _GEN_604; // @[Accumulator_Array.scala 57:76]
  assign io_isdone = acc_counter == 4'h8; // @[Accumulator_Array.scala 61:20]
  assign io_out_sum_0 = io_in_compute_done ? Acc_Result_0_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_1 = io_in_compute_done ? Acc_Result_0_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_2 = io_in_compute_done ? Acc_Result_0_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_3 = io_in_compute_done ? Acc_Result_0_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_4 = io_in_compute_done ? Acc_Result_0_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_5 = io_in_compute_done ? Acc_Result_0_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_6 = io_in_compute_done ? Acc_Result_0_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_7 = io_in_compute_done ? Acc_Result_0_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_8 = io_in_compute_done ? Acc_Result_1_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_9 = io_in_compute_done ? Acc_Result_1_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_10 = io_in_compute_done ? Acc_Result_1_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_11 = io_in_compute_done ? Acc_Result_1_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_12 = io_in_compute_done ? Acc_Result_1_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_13 = io_in_compute_done ? Acc_Result_1_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_14 = io_in_compute_done ? Acc_Result_1_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_15 = io_in_compute_done ? Acc_Result_1_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_16 = io_in_compute_done ? Acc_Result_2_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_17 = io_in_compute_done ? Acc_Result_2_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_18 = io_in_compute_done ? Acc_Result_2_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_19 = io_in_compute_done ? Acc_Result_2_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_20 = io_in_compute_done ? Acc_Result_2_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_21 = io_in_compute_done ? Acc_Result_2_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_22 = io_in_compute_done ? Acc_Result_2_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_23 = io_in_compute_done ? Acc_Result_2_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_24 = io_in_compute_done ? Acc_Result_3_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_25 = io_in_compute_done ? Acc_Result_3_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_26 = io_in_compute_done ? Acc_Result_3_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_27 = io_in_compute_done ? Acc_Result_3_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_28 = io_in_compute_done ? Acc_Result_3_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_29 = io_in_compute_done ? Acc_Result_3_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_30 = io_in_compute_done ? Acc_Result_3_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_31 = io_in_compute_done ? Acc_Result_3_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_32 = io_in_compute_done ? Acc_Result_4_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_33 = io_in_compute_done ? Acc_Result_4_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_34 = io_in_compute_done ? Acc_Result_4_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_35 = io_in_compute_done ? Acc_Result_4_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_36 = io_in_compute_done ? Acc_Result_4_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_37 = io_in_compute_done ? Acc_Result_4_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_38 = io_in_compute_done ? Acc_Result_4_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_39 = io_in_compute_done ? Acc_Result_4_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_40 = io_in_compute_done ? Acc_Result_5_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_41 = io_in_compute_done ? Acc_Result_5_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_42 = io_in_compute_done ? Acc_Result_5_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_43 = io_in_compute_done ? Acc_Result_5_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_44 = io_in_compute_done ? Acc_Result_5_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_45 = io_in_compute_done ? Acc_Result_5_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_46 = io_in_compute_done ? Acc_Result_5_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_47 = io_in_compute_done ? Acc_Result_5_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_48 = io_in_compute_done ? Acc_Result_6_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_49 = io_in_compute_done ? Acc_Result_6_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_50 = io_in_compute_done ? Acc_Result_6_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_51 = io_in_compute_done ? Acc_Result_6_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_52 = io_in_compute_done ? Acc_Result_6_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_53 = io_in_compute_done ? Acc_Result_6_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_54 = io_in_compute_done ? Acc_Result_6_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_55 = io_in_compute_done ? Acc_Result_6_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_56 = io_in_compute_done ? Acc_Result_7_0 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_57 = io_in_compute_done ? Acc_Result_7_1 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_58 = io_in_compute_done ? Acc_Result_7_2 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_59 = io_in_compute_done ? Acc_Result_7_3 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_60 = io_in_compute_done ? Acc_Result_7_4 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_61 = io_in_compute_done ? Acc_Result_7_5 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_62 = io_in_compute_done ? Acc_Result_7_6 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_out_sum_63 = io_in_compute_done ? Acc_Result_7_7 : 32'h0; // @[Accumulator_Array.scala 67:28 68:16 71:16]
  assign io_valid = io_in_compute_done; // @[Accumulator_Array.scala 67:28 69:14 72:14]
  always @(posedge clock) begin
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_0_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h0 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_0_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h0 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_0_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_0_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_1_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h1 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_1_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h1 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_1_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_1_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_2_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h2 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_2_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h2 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_2_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_2_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_3_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h3 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_3_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h3 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_3_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_3_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_4_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h4 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_4_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h4 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_4_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_4_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_5_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h5 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_5_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h5 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_5_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_5_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_0 <= Acc_Buffer_7_0; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_1 <= Acc_Buffer_7_1; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_2 <= Acc_Buffer_7_2; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_3 <= Acc_Buffer_7_3; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_4 <= Acc_Buffer_7_4; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_5 <= Acc_Buffer_7_5; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_6 <= Acc_Buffer_7_6; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_6_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h6 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_6_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h6 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_6_7 <= Acc_Buffer_7_7; // @[Accumulator_Array.scala 28:39]
      end else begin
        Acc_Buffer_6_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_0 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_0) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_0 <= io_in_psum_0; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_0[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_0[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_0 <= _GEN_22;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_1 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_1) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_1 <= io_in_psum_1; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_1[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_1[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_1 <= _GEN_54;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_2 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_2) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_2 <= io_in_psum_2; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_2[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_2[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_2 <= _GEN_86;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_3 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_3) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_3 <= io_in_psum_3; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_3[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_3[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_3 <= _GEN_118;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_4 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_4) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_4 <= io_in_psum_4; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_4[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_4[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_4 <= _GEN_150;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_5 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_5) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_5 <= io_in_psum_5; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_5[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_5[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_5 <= _GEN_182;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_6 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_6) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_6 <= io_in_psum_6; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_6[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_6[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_6 <= _GEN_214;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 20:27]
      Acc_Buffer_7_7 <= 16'h0; // @[Accumulator_Array.scala 20:27]
    end else if (io_in_valid_7) begin // @[Accumulator_Array.scala 25:26]
      if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 26:39]
        Acc_Buffer_7_7 <= io_in_psum_7; // @[Accumulator_Array.scala 26:39]
      end
    end else if (3'h7 == valid_counter_7[2:0]) begin // @[Accumulator_Array.scala 28:39]
      if (!(3'h7 == valid_counter_7[2:0])) begin // @[Accumulator_Array.scala 28:39]
        Acc_Buffer_7_7 <= _GEN_246;
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_0_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h0 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_0_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_1_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h1 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_1_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_2_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h2 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_2_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_3_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h3 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_3_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_4_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h4 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_4_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_5_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h5 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_5_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_6_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h6 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_6_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_0 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_0 <= _Acc_Result_0_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_1 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_1 <= _Acc_Result_1_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_2 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_2 <= _Acc_Result_2_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_3 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_3 <= _Acc_Result_3_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_4 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_4 <= _Acc_Result_4_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_5 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_5 <= _Acc_Result_5_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_6 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_6 <= _Acc_Result_6_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 21:27]
      Acc_Result_7_7 <= 32'h0; // @[Accumulator_Array.scala 21:27]
    end else if (_T_43) begin // @[Accumulator_Array.scala 55:29]
      if (3'h7 == _T_46[2:0]) begin // @[Accumulator_Array.scala 57:40]
        Acc_Result_7_7 <= _Acc_Result_7_T_7; // @[Accumulator_Array.scala 57:40]
      end
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_0 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_0 & valid_counter_0 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_0 <= _valid_counter_0_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_0 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_0 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_1 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_1 & valid_counter_1 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_1 <= _valid_counter_1_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_1 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_1 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_2 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_2 & valid_counter_2 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_2 <= _valid_counter_2_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_2 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_2 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_3 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_3 & valid_counter_3 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_3 <= _valid_counter_3_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_3 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_3 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_4 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_4 & valid_counter_4 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_4 <= _valid_counter_4_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_4 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_4 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_5 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_5 & valid_counter_5 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_5 <= _valid_counter_5_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_5 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_5 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_6 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_6 & valid_counter_6 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_6 <= _valid_counter_6_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_6 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_6 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 22:30]
      valid_counter_7 <= 4'h0; // @[Accumulator_Array.scala 22:30]
    end else if (io_in_valid_7 & valid_counter_7 < 4'h7) begin // @[Accumulator_Array.scala 34:67]
      valid_counter_7 <= _valid_counter_7_T_1; // @[Accumulator_Array.scala 35:24]
    end else if (valid_counter_7 == 4'h7) begin // @[Accumulator_Array.scala 36:55]
      valid_counter_7 <= 4'h0; // @[Accumulator_Array.scala 37:24]
    end
    if (reset) begin // @[Accumulator_Array.scala 43:28]
      acc_counter <= 4'h0; // @[Accumulator_Array.scala 43:28]
    end else if (io_in_acc & acc_counter == 4'h0) begin // @[Accumulator_Array.scala 45:44]
      acc_counter <= _acc_counter_T_1; // @[Accumulator_Array.scala 46:17]
    end else if (acc_counter == 4'h8) begin // @[Accumulator_Array.scala 47:43]
      acc_counter <= 4'h0; // @[Accumulator_Array.scala 48:17]
    end else if (acc_counter != 4'h0) begin // @[Accumulator_Array.scala 49:35]
      acc_counter <= _acc_counter_T_1; // @[Accumulator_Array.scala 50:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Acc_Buffer_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  Acc_Buffer_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  Acc_Buffer_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  Acc_Buffer_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  Acc_Buffer_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  Acc_Buffer_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  Acc_Buffer_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  Acc_Buffer_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  Acc_Buffer_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  Acc_Buffer_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  Acc_Buffer_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  Acc_Buffer_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  Acc_Buffer_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  Acc_Buffer_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  Acc_Buffer_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  Acc_Buffer_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  Acc_Buffer_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  Acc_Buffer_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  Acc_Buffer_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  Acc_Buffer_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  Acc_Buffer_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  Acc_Buffer_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  Acc_Buffer_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  Acc_Buffer_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  Acc_Buffer_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  Acc_Buffer_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  Acc_Buffer_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  Acc_Buffer_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  Acc_Buffer_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  Acc_Buffer_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  Acc_Buffer_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  Acc_Buffer_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  Acc_Buffer_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  Acc_Buffer_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  Acc_Buffer_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  Acc_Buffer_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  Acc_Buffer_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  Acc_Buffer_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  Acc_Buffer_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  Acc_Buffer_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  Acc_Buffer_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  Acc_Buffer_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  Acc_Buffer_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  Acc_Buffer_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  Acc_Buffer_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  Acc_Buffer_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  Acc_Buffer_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  Acc_Buffer_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  Acc_Buffer_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  Acc_Buffer_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  Acc_Buffer_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  Acc_Buffer_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  Acc_Buffer_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  Acc_Buffer_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  Acc_Buffer_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  Acc_Buffer_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  Acc_Buffer_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  Acc_Buffer_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  Acc_Buffer_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  Acc_Buffer_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  Acc_Buffer_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  Acc_Buffer_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  Acc_Buffer_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  Acc_Buffer_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  Acc_Result_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  Acc_Result_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  Acc_Result_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  Acc_Result_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  Acc_Result_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  Acc_Result_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  Acc_Result_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  Acc_Result_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  Acc_Result_1_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  Acc_Result_1_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  Acc_Result_1_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  Acc_Result_1_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  Acc_Result_1_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  Acc_Result_1_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  Acc_Result_1_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  Acc_Result_1_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  Acc_Result_2_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  Acc_Result_2_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  Acc_Result_2_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  Acc_Result_2_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  Acc_Result_2_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  Acc_Result_2_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  Acc_Result_2_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  Acc_Result_2_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  Acc_Result_3_0 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  Acc_Result_3_1 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  Acc_Result_3_2 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  Acc_Result_3_3 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  Acc_Result_3_4 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  Acc_Result_3_5 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  Acc_Result_3_6 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  Acc_Result_3_7 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  Acc_Result_4_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  Acc_Result_4_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  Acc_Result_4_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  Acc_Result_4_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  Acc_Result_4_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  Acc_Result_4_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  Acc_Result_4_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  Acc_Result_4_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  Acc_Result_5_0 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  Acc_Result_5_1 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  Acc_Result_5_2 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  Acc_Result_5_3 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  Acc_Result_5_4 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  Acc_Result_5_5 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  Acc_Result_5_6 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  Acc_Result_5_7 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  Acc_Result_6_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  Acc_Result_6_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  Acc_Result_6_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  Acc_Result_6_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  Acc_Result_6_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  Acc_Result_6_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  Acc_Result_6_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  Acc_Result_6_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  Acc_Result_7_0 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  Acc_Result_7_1 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  Acc_Result_7_2 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  Acc_Result_7_3 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  Acc_Result_7_4 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  Acc_Result_7_5 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  Acc_Result_7_6 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  Acc_Result_7_7 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_counter_0 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  valid_counter_1 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  valid_counter_2 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  valid_counter_3 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  valid_counter_4 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  valid_counter_5 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  valid_counter_6 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  valid_counter_7 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  acc_counter = _RAND_136[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mini_TPU(
  input         clock,
  input         reset,
  input         io_Compute,
  output        io_Data_x_ready,
  input         io_Data_x_valid,
  input  [7:0]  io_Data_x_bits_0,
  input  [7:0]  io_Data_x_bits_1,
  input  [7:0]  io_Data_x_bits_2,
  input  [7:0]  io_Data_x_bits_3,
  input  [7:0]  io_Data_x_bits_4,
  input  [7:0]  io_Data_x_bits_5,
  input  [7:0]  io_Data_x_bits_6,
  input  [7:0]  io_Data_x_bits_7,
  input  [7:0]  io_Data_x_bits_8,
  input  [7:0]  io_Data_x_bits_9,
  input  [7:0]  io_Data_x_bits_10,
  input  [7:0]  io_Data_x_bits_11,
  input  [7:0]  io_Data_x_bits_12,
  input  [7:0]  io_Data_x_bits_13,
  input  [7:0]  io_Data_x_bits_14,
  input  [7:0]  io_Data_x_bits_15,
  input  [7:0]  io_Data_x_bits_16,
  input  [7:0]  io_Data_x_bits_17,
  input  [7:0]  io_Data_x_bits_18,
  input  [7:0]  io_Data_x_bits_19,
  input  [7:0]  io_Data_x_bits_20,
  input  [7:0]  io_Data_x_bits_21,
  input  [7:0]  io_Data_x_bits_22,
  input  [7:0]  io_Data_x_bits_23,
  input  [7:0]  io_Data_x_bits_24,
  input  [7:0]  io_Data_x_bits_25,
  input  [7:0]  io_Data_x_bits_26,
  input  [7:0]  io_Data_x_bits_27,
  input  [7:0]  io_Data_x_bits_28,
  input  [7:0]  io_Data_x_bits_29,
  input  [7:0]  io_Data_x_bits_30,
  input  [7:0]  io_Data_x_bits_31,
  input  [7:0]  io_Data_x_bits_32,
  input  [7:0]  io_Data_x_bits_33,
  input  [7:0]  io_Data_x_bits_34,
  input  [7:0]  io_Data_x_bits_35,
  input  [7:0]  io_Data_x_bits_36,
  input  [7:0]  io_Data_x_bits_37,
  input  [7:0]  io_Data_x_bits_38,
  input  [7:0]  io_Data_x_bits_39,
  input  [7:0]  io_Data_x_bits_40,
  input  [7:0]  io_Data_x_bits_41,
  input  [7:0]  io_Data_x_bits_42,
  input  [7:0]  io_Data_x_bits_43,
  input  [7:0]  io_Data_x_bits_44,
  input  [7:0]  io_Data_x_bits_45,
  input  [7:0]  io_Data_x_bits_46,
  input  [7:0]  io_Data_x_bits_47,
  input  [7:0]  io_Data_x_bits_48,
  input  [7:0]  io_Data_x_bits_49,
  input  [7:0]  io_Data_x_bits_50,
  input  [7:0]  io_Data_x_bits_51,
  input  [7:0]  io_Data_x_bits_52,
  input  [7:0]  io_Data_x_bits_53,
  input  [7:0]  io_Data_x_bits_54,
  input  [7:0]  io_Data_x_bits_55,
  input  [7:0]  io_Data_x_bits_56,
  input  [7:0]  io_Data_x_bits_57,
  input  [7:0]  io_Data_x_bits_58,
  input  [7:0]  io_Data_x_bits_59,
  input  [7:0]  io_Data_x_bits_60,
  input  [7:0]  io_Data_x_bits_61,
  input  [7:0]  io_Data_x_bits_62,
  input  [7:0]  io_Data_x_bits_63,
  output        io_Weight_x_ready,
  input         io_Weight_x_valid,
  input  [7:0]  io_Weight_x_bits_0,
  input  [7:0]  io_Weight_x_bits_1,
  input  [7:0]  io_Weight_x_bits_2,
  input  [7:0]  io_Weight_x_bits_3,
  input  [7:0]  io_Weight_x_bits_4,
  input  [7:0]  io_Weight_x_bits_5,
  input  [7:0]  io_Weight_x_bits_6,
  input  [7:0]  io_Weight_x_bits_7,
  input  [7:0]  io_Weight_x_bits_8,
  input  [7:0]  io_Weight_x_bits_9,
  input  [7:0]  io_Weight_x_bits_10,
  input  [7:0]  io_Weight_x_bits_11,
  input  [7:0]  io_Weight_x_bits_12,
  input  [7:0]  io_Weight_x_bits_13,
  input  [7:0]  io_Weight_x_bits_14,
  input  [7:0]  io_Weight_x_bits_15,
  input  [7:0]  io_Weight_x_bits_16,
  input  [7:0]  io_Weight_x_bits_17,
  input  [7:0]  io_Weight_x_bits_18,
  input  [7:0]  io_Weight_x_bits_19,
  input  [7:0]  io_Weight_x_bits_20,
  input  [7:0]  io_Weight_x_bits_21,
  input  [7:0]  io_Weight_x_bits_22,
  input  [7:0]  io_Weight_x_bits_23,
  input  [7:0]  io_Weight_x_bits_24,
  input  [7:0]  io_Weight_x_bits_25,
  input  [7:0]  io_Weight_x_bits_26,
  input  [7:0]  io_Weight_x_bits_27,
  input  [7:0]  io_Weight_x_bits_28,
  input  [7:0]  io_Weight_x_bits_29,
  input  [7:0]  io_Weight_x_bits_30,
  input  [7:0]  io_Weight_x_bits_31,
  input  [7:0]  io_Weight_x_bits_32,
  input  [7:0]  io_Weight_x_bits_33,
  input  [7:0]  io_Weight_x_bits_34,
  input  [7:0]  io_Weight_x_bits_35,
  input  [7:0]  io_Weight_x_bits_36,
  input  [7:0]  io_Weight_x_bits_37,
  input  [7:0]  io_Weight_x_bits_38,
  input  [7:0]  io_Weight_x_bits_39,
  input  [7:0]  io_Weight_x_bits_40,
  input  [7:0]  io_Weight_x_bits_41,
  input  [7:0]  io_Weight_x_bits_42,
  input  [7:0]  io_Weight_x_bits_43,
  input  [7:0]  io_Weight_x_bits_44,
  input  [7:0]  io_Weight_x_bits_45,
  input  [7:0]  io_Weight_x_bits_46,
  input  [7:0]  io_Weight_x_bits_47,
  input  [7:0]  io_Weight_x_bits_48,
  input  [7:0]  io_Weight_x_bits_49,
  input  [7:0]  io_Weight_x_bits_50,
  input  [7:0]  io_Weight_x_bits_51,
  input  [7:0]  io_Weight_x_bits_52,
  input  [7:0]  io_Weight_x_bits_53,
  input  [7:0]  io_Weight_x_bits_54,
  input  [7:0]  io_Weight_x_bits_55,
  input  [7:0]  io_Weight_x_bits_56,
  input  [7:0]  io_Weight_x_bits_57,
  input  [7:0]  io_Weight_x_bits_58,
  input  [7:0]  io_Weight_x_bits_59,
  input  [7:0]  io_Weight_x_bits_60,
  input  [7:0]  io_Weight_x_bits_61,
  input  [7:0]  io_Weight_x_bits_62,
  input  [7:0]  io_Weight_x_bits_63,
  input         io_Sum_x_ready,
  output        io_Sum_x_valid,
  output [31:0] io_Sum_x_bits_0,
  output [31:0] io_Sum_x_bits_1,
  output [31:0] io_Sum_x_bits_2,
  output [31:0] io_Sum_x_bits_3,
  output [31:0] io_Sum_x_bits_4,
  output [31:0] io_Sum_x_bits_5,
  output [31:0] io_Sum_x_bits_6,
  output [31:0] io_Sum_x_bits_7,
  output [31:0] io_Sum_x_bits_8,
  output [31:0] io_Sum_x_bits_9,
  output [31:0] io_Sum_x_bits_10,
  output [31:0] io_Sum_x_bits_11,
  output [31:0] io_Sum_x_bits_12,
  output [31:0] io_Sum_x_bits_13,
  output [31:0] io_Sum_x_bits_14,
  output [31:0] io_Sum_x_bits_15,
  output [31:0] io_Sum_x_bits_16,
  output [31:0] io_Sum_x_bits_17,
  output [31:0] io_Sum_x_bits_18,
  output [31:0] io_Sum_x_bits_19,
  output [31:0] io_Sum_x_bits_20,
  output [31:0] io_Sum_x_bits_21,
  output [31:0] io_Sum_x_bits_22,
  output [31:0] io_Sum_x_bits_23,
  output [31:0] io_Sum_x_bits_24,
  output [31:0] io_Sum_x_bits_25,
  output [31:0] io_Sum_x_bits_26,
  output [31:0] io_Sum_x_bits_27,
  output [31:0] io_Sum_x_bits_28,
  output [31:0] io_Sum_x_bits_29,
  output [31:0] io_Sum_x_bits_30,
  output [31:0] io_Sum_x_bits_31,
  output [31:0] io_Sum_x_bits_32,
  output [31:0] io_Sum_x_bits_33,
  output [31:0] io_Sum_x_bits_34,
  output [31:0] io_Sum_x_bits_35,
  output [31:0] io_Sum_x_bits_36,
  output [31:0] io_Sum_x_bits_37,
  output [31:0] io_Sum_x_bits_38,
  output [31:0] io_Sum_x_bits_39,
  output [31:0] io_Sum_x_bits_40,
  output [31:0] io_Sum_x_bits_41,
  output [31:0] io_Sum_x_bits_42,
  output [31:0] io_Sum_x_bits_43,
  output [31:0] io_Sum_x_bits_44,
  output [31:0] io_Sum_x_bits_45,
  output [31:0] io_Sum_x_bits_46,
  output [31:0] io_Sum_x_bits_47,
  output [31:0] io_Sum_x_bits_48,
  output [31:0] io_Sum_x_bits_49,
  output [31:0] io_Sum_x_bits_50,
  output [31:0] io_Sum_x_bits_51,
  output [31:0] io_Sum_x_bits_52,
  output [31:0] io_Sum_x_bits_53,
  output [31:0] io_Sum_x_bits_54,
  output [31:0] io_Sum_x_bits_55,
  output [31:0] io_Sum_x_bits_56,
  output [31:0] io_Sum_x_bits_57,
  output [31:0] io_Sum_x_bits_58,
  output [31:0] io_Sum_x_bits_59,
  output [31:0] io_Sum_x_bits_60,
  output [31:0] io_Sum_x_bits_61,
  output [31:0] io_Sum_x_bits_62,
  output [31:0] io_Sum_x_bits_63
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  activation_buffer_clock; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_reset; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_wen; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_ren; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_0; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_1; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_2; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_3; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_4; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_5; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_6; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_7; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_8; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_9; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_10; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_11; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_12; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_13; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_14; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_15; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_16; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_17; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_18; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_19; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_20; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_21; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_22; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_23; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_24; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_25; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_26; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_27; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_28; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_29; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_30; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_31; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_32; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_33; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_34; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_35; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_36; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_37; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_38; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_39; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_40; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_41; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_42; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_43; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_44; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_45; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_46; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_47; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_48; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_49; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_50; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_51; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_52; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_53; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_54; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_55; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_56; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_57; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_58; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_59; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_60; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_61; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_62; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_in_data_x_63; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_0; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_1; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_2; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_3; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_4; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_5; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_6; // @[Mini_TPU.scala 17:33]
  wire [7:0] activation_buffer_io_out_activate_7; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_out_flow; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_isfull; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_isempty; // @[Mini_TPU.scala 17:33]
  wire  activation_buffer_io_isdone; // @[Mini_TPU.scala 17:33]
  wire  weight_buffer_clock; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_reset; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_wen; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_ren; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_0; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_1; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_2; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_3; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_4; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_5; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_6; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_7; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_8; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_9; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_10; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_11; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_12; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_13; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_14; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_15; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_16; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_17; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_18; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_19; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_20; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_21; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_22; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_23; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_24; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_25; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_26; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_27; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_28; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_29; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_30; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_31; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_32; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_33; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_34; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_35; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_36; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_37; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_38; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_39; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_40; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_41; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_42; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_43; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_44; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_45; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_46; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_47; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_48; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_49; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_50; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_51; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_52; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_53; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_54; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_55; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_56; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_57; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_58; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_59; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_60; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_61; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_62; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_in_weight_x_63; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_0; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_1; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_2; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_3; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_4; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_5; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_6; // @[Mini_TPU.scala 18:29]
  wire [7:0] weight_buffer_io_out_weight_7; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_out_shift; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_isfull; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_isempty; // @[Mini_TPU.scala 18:29]
  wire  weight_buffer_io_isdone; // @[Mini_TPU.scala 18:29]
  wire  systolic_array_clock; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_reset; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_0; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_1; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_2; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_3; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_4; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_5; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_6; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_activate_7; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_0; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_1; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_2; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_3; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_4; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_5; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_6; // @[Mini_TPU.scala 19:30]
  wire [7:0] systolic_array_io_weight_7; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_flow; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_shift; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_0; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_1; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_2; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_3; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_4; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_5; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_6; // @[Mini_TPU.scala 19:30]
  wire [15:0] systolic_array_io_psum_7; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_0; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_1; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_2; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_3; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_4; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_5; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_6; // @[Mini_TPU.scala 19:30]
  wire  systolic_array_io_valid_7; // @[Mini_TPU.scala 19:30]
  wire  accumulation_array_clock; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_reset; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_0; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_1; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_2; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_3; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_4; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_5; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_6; // @[Mini_TPU.scala 20:34]
  wire [15:0] accumulation_array_io_in_psum_7; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_0; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_1; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_2; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_3; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_4; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_5; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_6; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_valid_7; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_acc; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_in_compute_done; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_isdone; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_0; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_1; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_2; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_3; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_4; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_5; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_6; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_7; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_8; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_9; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_10; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_11; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_12; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_13; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_14; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_15; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_16; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_17; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_18; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_19; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_20; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_21; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_22; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_23; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_24; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_25; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_26; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_27; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_28; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_29; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_30; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_31; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_32; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_33; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_34; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_35; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_36; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_37; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_38; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_39; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_40; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_41; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_42; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_43; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_44; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_45; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_46; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_47; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_48; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_49; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_50; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_51; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_52; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_53; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_54; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_55; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_56; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_57; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_58; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_59; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_60; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_61; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_62; // @[Mini_TPU.scala 20:34]
  wire [31:0] accumulation_array_io_out_sum_63; // @[Mini_TPU.scala 20:34]
  wire  accumulation_array_io_valid; // @[Mini_TPU.scala 20:34]
  reg [2:0] stateReg; // @[Mini_TPU.scala 24:25]
  wire  _T_1 = ~activation_buffer_io_isempty; // @[Mini_TPU.scala 35:27]
  wire  _T_3 = ~weight_buffer_io_isempty; // @[Mini_TPU.scala 35:62]
  wire  _T_4 = io_Compute & ~activation_buffer_io_isempty & ~weight_buffer_io_isempty; // @[Mini_TPU.scala 35:58]
  wire  _GEN_2 = weight_buffer_io_isdone; // @[Mini_TPU.scala 27:28 44:37 45:34]
  wire  _GEN_4 = activation_buffer_io_isdone; // @[Mini_TPU.scala 29:32 53:41 54:38]
  wire [2:0] _GEN_5 = activation_buffer_io_isdone ? 3'h3 : 3'h2; // @[Mini_TPU.scala 53:41 55:18 57:18]
  wire  _T_10 = _T_1 & _T_3; // @[Mini_TPU.scala 63:46]
  wire [2:0] _GEN_7 = _T_1 & _T_3 ? 3'h1 : 3'h4; // @[Mini_TPU.scala 63:78 65:20 67:20]
  wire  _GEN_8 = accumulation_array_io_isdone & _T_10; // @[Mini_TPU.scala 28:24 62:42]
  wire [2:0] _GEN_9 = accumulation_array_io_isdone ? _GEN_7 : 3'h3; // @[Mini_TPU.scala 62:42 70:18]
  wire [2:0] _GEN_11 = 3'h4 == stateReg ? 3'h0 : stateReg; // @[Mini_TPU.scala 32:20 75:16 24:25]
  wire [2:0] _GEN_14 = 3'h3 == stateReg ? _GEN_9 : _GEN_11; // @[Mini_TPU.scala 32:20]
  wire  _GEN_15 = 3'h3 == stateReg ? 1'h0 : 3'h4 == stateReg; // @[Mini_TPU.scala 32:20 30:41]
  wire  _GEN_19 = 3'h2 == stateReg ? 1'h0 : 3'h3 == stateReg & _GEN_8; // @[Mini_TPU.scala 32:20 28:24]
  wire  _GEN_20 = 3'h2 == stateReg ? 1'h0 : _GEN_15; // @[Mini_TPU.scala 32:20 30:41]
  wire  _GEN_21 = 3'h1 == stateReg ? 1'h0 : _GEN_19; // @[Mini_TPU.scala 32:20 43:28]
  wire  _GEN_24 = 3'h1 == stateReg ? 1'h0 : 3'h2 == stateReg & _GEN_4; // @[Mini_TPU.scala 32:20 29:32]
  wire  _GEN_25 = 3'h1 == stateReg ? 1'h0 : _GEN_20; // @[Mini_TPU.scala 32:20 30:41]
  wire  _T_12 = io_Sum_x_ready & io_Sum_x_valid; // @[Decoupled.scala 52:35]
  Activation_Buffer activation_buffer ( // @[Mini_TPU.scala 17:33]
    .clock(activation_buffer_clock),
    .reset(activation_buffer_reset),
    .io_wen(activation_buffer_io_wen),
    .io_ren(activation_buffer_io_ren),
    .io_in_data_x_0(activation_buffer_io_in_data_x_0),
    .io_in_data_x_1(activation_buffer_io_in_data_x_1),
    .io_in_data_x_2(activation_buffer_io_in_data_x_2),
    .io_in_data_x_3(activation_buffer_io_in_data_x_3),
    .io_in_data_x_4(activation_buffer_io_in_data_x_4),
    .io_in_data_x_5(activation_buffer_io_in_data_x_5),
    .io_in_data_x_6(activation_buffer_io_in_data_x_6),
    .io_in_data_x_7(activation_buffer_io_in_data_x_7),
    .io_in_data_x_8(activation_buffer_io_in_data_x_8),
    .io_in_data_x_9(activation_buffer_io_in_data_x_9),
    .io_in_data_x_10(activation_buffer_io_in_data_x_10),
    .io_in_data_x_11(activation_buffer_io_in_data_x_11),
    .io_in_data_x_12(activation_buffer_io_in_data_x_12),
    .io_in_data_x_13(activation_buffer_io_in_data_x_13),
    .io_in_data_x_14(activation_buffer_io_in_data_x_14),
    .io_in_data_x_15(activation_buffer_io_in_data_x_15),
    .io_in_data_x_16(activation_buffer_io_in_data_x_16),
    .io_in_data_x_17(activation_buffer_io_in_data_x_17),
    .io_in_data_x_18(activation_buffer_io_in_data_x_18),
    .io_in_data_x_19(activation_buffer_io_in_data_x_19),
    .io_in_data_x_20(activation_buffer_io_in_data_x_20),
    .io_in_data_x_21(activation_buffer_io_in_data_x_21),
    .io_in_data_x_22(activation_buffer_io_in_data_x_22),
    .io_in_data_x_23(activation_buffer_io_in_data_x_23),
    .io_in_data_x_24(activation_buffer_io_in_data_x_24),
    .io_in_data_x_25(activation_buffer_io_in_data_x_25),
    .io_in_data_x_26(activation_buffer_io_in_data_x_26),
    .io_in_data_x_27(activation_buffer_io_in_data_x_27),
    .io_in_data_x_28(activation_buffer_io_in_data_x_28),
    .io_in_data_x_29(activation_buffer_io_in_data_x_29),
    .io_in_data_x_30(activation_buffer_io_in_data_x_30),
    .io_in_data_x_31(activation_buffer_io_in_data_x_31),
    .io_in_data_x_32(activation_buffer_io_in_data_x_32),
    .io_in_data_x_33(activation_buffer_io_in_data_x_33),
    .io_in_data_x_34(activation_buffer_io_in_data_x_34),
    .io_in_data_x_35(activation_buffer_io_in_data_x_35),
    .io_in_data_x_36(activation_buffer_io_in_data_x_36),
    .io_in_data_x_37(activation_buffer_io_in_data_x_37),
    .io_in_data_x_38(activation_buffer_io_in_data_x_38),
    .io_in_data_x_39(activation_buffer_io_in_data_x_39),
    .io_in_data_x_40(activation_buffer_io_in_data_x_40),
    .io_in_data_x_41(activation_buffer_io_in_data_x_41),
    .io_in_data_x_42(activation_buffer_io_in_data_x_42),
    .io_in_data_x_43(activation_buffer_io_in_data_x_43),
    .io_in_data_x_44(activation_buffer_io_in_data_x_44),
    .io_in_data_x_45(activation_buffer_io_in_data_x_45),
    .io_in_data_x_46(activation_buffer_io_in_data_x_46),
    .io_in_data_x_47(activation_buffer_io_in_data_x_47),
    .io_in_data_x_48(activation_buffer_io_in_data_x_48),
    .io_in_data_x_49(activation_buffer_io_in_data_x_49),
    .io_in_data_x_50(activation_buffer_io_in_data_x_50),
    .io_in_data_x_51(activation_buffer_io_in_data_x_51),
    .io_in_data_x_52(activation_buffer_io_in_data_x_52),
    .io_in_data_x_53(activation_buffer_io_in_data_x_53),
    .io_in_data_x_54(activation_buffer_io_in_data_x_54),
    .io_in_data_x_55(activation_buffer_io_in_data_x_55),
    .io_in_data_x_56(activation_buffer_io_in_data_x_56),
    .io_in_data_x_57(activation_buffer_io_in_data_x_57),
    .io_in_data_x_58(activation_buffer_io_in_data_x_58),
    .io_in_data_x_59(activation_buffer_io_in_data_x_59),
    .io_in_data_x_60(activation_buffer_io_in_data_x_60),
    .io_in_data_x_61(activation_buffer_io_in_data_x_61),
    .io_in_data_x_62(activation_buffer_io_in_data_x_62),
    .io_in_data_x_63(activation_buffer_io_in_data_x_63),
    .io_out_activate_0(activation_buffer_io_out_activate_0),
    .io_out_activate_1(activation_buffer_io_out_activate_1),
    .io_out_activate_2(activation_buffer_io_out_activate_2),
    .io_out_activate_3(activation_buffer_io_out_activate_3),
    .io_out_activate_4(activation_buffer_io_out_activate_4),
    .io_out_activate_5(activation_buffer_io_out_activate_5),
    .io_out_activate_6(activation_buffer_io_out_activate_6),
    .io_out_activate_7(activation_buffer_io_out_activate_7),
    .io_out_flow(activation_buffer_io_out_flow),
    .io_isfull(activation_buffer_io_isfull),
    .io_isempty(activation_buffer_io_isempty),
    .io_isdone(activation_buffer_io_isdone)
  );
  Weight_Buffer weight_buffer ( // @[Mini_TPU.scala 18:29]
    .clock(weight_buffer_clock),
    .reset(weight_buffer_reset),
    .io_wen(weight_buffer_io_wen),
    .io_ren(weight_buffer_io_ren),
    .io_in_weight_x_0(weight_buffer_io_in_weight_x_0),
    .io_in_weight_x_1(weight_buffer_io_in_weight_x_1),
    .io_in_weight_x_2(weight_buffer_io_in_weight_x_2),
    .io_in_weight_x_3(weight_buffer_io_in_weight_x_3),
    .io_in_weight_x_4(weight_buffer_io_in_weight_x_4),
    .io_in_weight_x_5(weight_buffer_io_in_weight_x_5),
    .io_in_weight_x_6(weight_buffer_io_in_weight_x_6),
    .io_in_weight_x_7(weight_buffer_io_in_weight_x_7),
    .io_in_weight_x_8(weight_buffer_io_in_weight_x_8),
    .io_in_weight_x_9(weight_buffer_io_in_weight_x_9),
    .io_in_weight_x_10(weight_buffer_io_in_weight_x_10),
    .io_in_weight_x_11(weight_buffer_io_in_weight_x_11),
    .io_in_weight_x_12(weight_buffer_io_in_weight_x_12),
    .io_in_weight_x_13(weight_buffer_io_in_weight_x_13),
    .io_in_weight_x_14(weight_buffer_io_in_weight_x_14),
    .io_in_weight_x_15(weight_buffer_io_in_weight_x_15),
    .io_in_weight_x_16(weight_buffer_io_in_weight_x_16),
    .io_in_weight_x_17(weight_buffer_io_in_weight_x_17),
    .io_in_weight_x_18(weight_buffer_io_in_weight_x_18),
    .io_in_weight_x_19(weight_buffer_io_in_weight_x_19),
    .io_in_weight_x_20(weight_buffer_io_in_weight_x_20),
    .io_in_weight_x_21(weight_buffer_io_in_weight_x_21),
    .io_in_weight_x_22(weight_buffer_io_in_weight_x_22),
    .io_in_weight_x_23(weight_buffer_io_in_weight_x_23),
    .io_in_weight_x_24(weight_buffer_io_in_weight_x_24),
    .io_in_weight_x_25(weight_buffer_io_in_weight_x_25),
    .io_in_weight_x_26(weight_buffer_io_in_weight_x_26),
    .io_in_weight_x_27(weight_buffer_io_in_weight_x_27),
    .io_in_weight_x_28(weight_buffer_io_in_weight_x_28),
    .io_in_weight_x_29(weight_buffer_io_in_weight_x_29),
    .io_in_weight_x_30(weight_buffer_io_in_weight_x_30),
    .io_in_weight_x_31(weight_buffer_io_in_weight_x_31),
    .io_in_weight_x_32(weight_buffer_io_in_weight_x_32),
    .io_in_weight_x_33(weight_buffer_io_in_weight_x_33),
    .io_in_weight_x_34(weight_buffer_io_in_weight_x_34),
    .io_in_weight_x_35(weight_buffer_io_in_weight_x_35),
    .io_in_weight_x_36(weight_buffer_io_in_weight_x_36),
    .io_in_weight_x_37(weight_buffer_io_in_weight_x_37),
    .io_in_weight_x_38(weight_buffer_io_in_weight_x_38),
    .io_in_weight_x_39(weight_buffer_io_in_weight_x_39),
    .io_in_weight_x_40(weight_buffer_io_in_weight_x_40),
    .io_in_weight_x_41(weight_buffer_io_in_weight_x_41),
    .io_in_weight_x_42(weight_buffer_io_in_weight_x_42),
    .io_in_weight_x_43(weight_buffer_io_in_weight_x_43),
    .io_in_weight_x_44(weight_buffer_io_in_weight_x_44),
    .io_in_weight_x_45(weight_buffer_io_in_weight_x_45),
    .io_in_weight_x_46(weight_buffer_io_in_weight_x_46),
    .io_in_weight_x_47(weight_buffer_io_in_weight_x_47),
    .io_in_weight_x_48(weight_buffer_io_in_weight_x_48),
    .io_in_weight_x_49(weight_buffer_io_in_weight_x_49),
    .io_in_weight_x_50(weight_buffer_io_in_weight_x_50),
    .io_in_weight_x_51(weight_buffer_io_in_weight_x_51),
    .io_in_weight_x_52(weight_buffer_io_in_weight_x_52),
    .io_in_weight_x_53(weight_buffer_io_in_weight_x_53),
    .io_in_weight_x_54(weight_buffer_io_in_weight_x_54),
    .io_in_weight_x_55(weight_buffer_io_in_weight_x_55),
    .io_in_weight_x_56(weight_buffer_io_in_weight_x_56),
    .io_in_weight_x_57(weight_buffer_io_in_weight_x_57),
    .io_in_weight_x_58(weight_buffer_io_in_weight_x_58),
    .io_in_weight_x_59(weight_buffer_io_in_weight_x_59),
    .io_in_weight_x_60(weight_buffer_io_in_weight_x_60),
    .io_in_weight_x_61(weight_buffer_io_in_weight_x_61),
    .io_in_weight_x_62(weight_buffer_io_in_weight_x_62),
    .io_in_weight_x_63(weight_buffer_io_in_weight_x_63),
    .io_out_weight_0(weight_buffer_io_out_weight_0),
    .io_out_weight_1(weight_buffer_io_out_weight_1),
    .io_out_weight_2(weight_buffer_io_out_weight_2),
    .io_out_weight_3(weight_buffer_io_out_weight_3),
    .io_out_weight_4(weight_buffer_io_out_weight_4),
    .io_out_weight_5(weight_buffer_io_out_weight_5),
    .io_out_weight_6(weight_buffer_io_out_weight_6),
    .io_out_weight_7(weight_buffer_io_out_weight_7),
    .io_out_shift(weight_buffer_io_out_shift),
    .io_isfull(weight_buffer_io_isfull),
    .io_isempty(weight_buffer_io_isempty),
    .io_isdone(weight_buffer_io_isdone)
  );
  Systolic_Array systolic_array ( // @[Mini_TPU.scala 19:30]
    .clock(systolic_array_clock),
    .reset(systolic_array_reset),
    .io_activate_0(systolic_array_io_activate_0),
    .io_activate_1(systolic_array_io_activate_1),
    .io_activate_2(systolic_array_io_activate_2),
    .io_activate_3(systolic_array_io_activate_3),
    .io_activate_4(systolic_array_io_activate_4),
    .io_activate_5(systolic_array_io_activate_5),
    .io_activate_6(systolic_array_io_activate_6),
    .io_activate_7(systolic_array_io_activate_7),
    .io_weight_0(systolic_array_io_weight_0),
    .io_weight_1(systolic_array_io_weight_1),
    .io_weight_2(systolic_array_io_weight_2),
    .io_weight_3(systolic_array_io_weight_3),
    .io_weight_4(systolic_array_io_weight_4),
    .io_weight_5(systolic_array_io_weight_5),
    .io_weight_6(systolic_array_io_weight_6),
    .io_weight_7(systolic_array_io_weight_7),
    .io_flow(systolic_array_io_flow),
    .io_shift(systolic_array_io_shift),
    .io_psum_0(systolic_array_io_psum_0),
    .io_psum_1(systolic_array_io_psum_1),
    .io_psum_2(systolic_array_io_psum_2),
    .io_psum_3(systolic_array_io_psum_3),
    .io_psum_4(systolic_array_io_psum_4),
    .io_psum_5(systolic_array_io_psum_5),
    .io_psum_6(systolic_array_io_psum_6),
    .io_psum_7(systolic_array_io_psum_7),
    .io_valid_0(systolic_array_io_valid_0),
    .io_valid_1(systolic_array_io_valid_1),
    .io_valid_2(systolic_array_io_valid_2),
    .io_valid_3(systolic_array_io_valid_3),
    .io_valid_4(systolic_array_io_valid_4),
    .io_valid_5(systolic_array_io_valid_5),
    .io_valid_6(systolic_array_io_valid_6),
    .io_valid_7(systolic_array_io_valid_7)
  );
  Accumulator_Array accumulation_array ( // @[Mini_TPU.scala 20:34]
    .clock(accumulation_array_clock),
    .reset(accumulation_array_reset),
    .io_in_psum_0(accumulation_array_io_in_psum_0),
    .io_in_psum_1(accumulation_array_io_in_psum_1),
    .io_in_psum_2(accumulation_array_io_in_psum_2),
    .io_in_psum_3(accumulation_array_io_in_psum_3),
    .io_in_psum_4(accumulation_array_io_in_psum_4),
    .io_in_psum_5(accumulation_array_io_in_psum_5),
    .io_in_psum_6(accumulation_array_io_in_psum_6),
    .io_in_psum_7(accumulation_array_io_in_psum_7),
    .io_in_valid_0(accumulation_array_io_in_valid_0),
    .io_in_valid_1(accumulation_array_io_in_valid_1),
    .io_in_valid_2(accumulation_array_io_in_valid_2),
    .io_in_valid_3(accumulation_array_io_in_valid_3),
    .io_in_valid_4(accumulation_array_io_in_valid_4),
    .io_in_valid_5(accumulation_array_io_in_valid_5),
    .io_in_valid_6(accumulation_array_io_in_valid_6),
    .io_in_valid_7(accumulation_array_io_in_valid_7),
    .io_in_acc(accumulation_array_io_in_acc),
    .io_in_compute_done(accumulation_array_io_in_compute_done),
    .io_isdone(accumulation_array_io_isdone),
    .io_out_sum_0(accumulation_array_io_out_sum_0),
    .io_out_sum_1(accumulation_array_io_out_sum_1),
    .io_out_sum_2(accumulation_array_io_out_sum_2),
    .io_out_sum_3(accumulation_array_io_out_sum_3),
    .io_out_sum_4(accumulation_array_io_out_sum_4),
    .io_out_sum_5(accumulation_array_io_out_sum_5),
    .io_out_sum_6(accumulation_array_io_out_sum_6),
    .io_out_sum_7(accumulation_array_io_out_sum_7),
    .io_out_sum_8(accumulation_array_io_out_sum_8),
    .io_out_sum_9(accumulation_array_io_out_sum_9),
    .io_out_sum_10(accumulation_array_io_out_sum_10),
    .io_out_sum_11(accumulation_array_io_out_sum_11),
    .io_out_sum_12(accumulation_array_io_out_sum_12),
    .io_out_sum_13(accumulation_array_io_out_sum_13),
    .io_out_sum_14(accumulation_array_io_out_sum_14),
    .io_out_sum_15(accumulation_array_io_out_sum_15),
    .io_out_sum_16(accumulation_array_io_out_sum_16),
    .io_out_sum_17(accumulation_array_io_out_sum_17),
    .io_out_sum_18(accumulation_array_io_out_sum_18),
    .io_out_sum_19(accumulation_array_io_out_sum_19),
    .io_out_sum_20(accumulation_array_io_out_sum_20),
    .io_out_sum_21(accumulation_array_io_out_sum_21),
    .io_out_sum_22(accumulation_array_io_out_sum_22),
    .io_out_sum_23(accumulation_array_io_out_sum_23),
    .io_out_sum_24(accumulation_array_io_out_sum_24),
    .io_out_sum_25(accumulation_array_io_out_sum_25),
    .io_out_sum_26(accumulation_array_io_out_sum_26),
    .io_out_sum_27(accumulation_array_io_out_sum_27),
    .io_out_sum_28(accumulation_array_io_out_sum_28),
    .io_out_sum_29(accumulation_array_io_out_sum_29),
    .io_out_sum_30(accumulation_array_io_out_sum_30),
    .io_out_sum_31(accumulation_array_io_out_sum_31),
    .io_out_sum_32(accumulation_array_io_out_sum_32),
    .io_out_sum_33(accumulation_array_io_out_sum_33),
    .io_out_sum_34(accumulation_array_io_out_sum_34),
    .io_out_sum_35(accumulation_array_io_out_sum_35),
    .io_out_sum_36(accumulation_array_io_out_sum_36),
    .io_out_sum_37(accumulation_array_io_out_sum_37),
    .io_out_sum_38(accumulation_array_io_out_sum_38),
    .io_out_sum_39(accumulation_array_io_out_sum_39),
    .io_out_sum_40(accumulation_array_io_out_sum_40),
    .io_out_sum_41(accumulation_array_io_out_sum_41),
    .io_out_sum_42(accumulation_array_io_out_sum_42),
    .io_out_sum_43(accumulation_array_io_out_sum_43),
    .io_out_sum_44(accumulation_array_io_out_sum_44),
    .io_out_sum_45(accumulation_array_io_out_sum_45),
    .io_out_sum_46(accumulation_array_io_out_sum_46),
    .io_out_sum_47(accumulation_array_io_out_sum_47),
    .io_out_sum_48(accumulation_array_io_out_sum_48),
    .io_out_sum_49(accumulation_array_io_out_sum_49),
    .io_out_sum_50(accumulation_array_io_out_sum_50),
    .io_out_sum_51(accumulation_array_io_out_sum_51),
    .io_out_sum_52(accumulation_array_io_out_sum_52),
    .io_out_sum_53(accumulation_array_io_out_sum_53),
    .io_out_sum_54(accumulation_array_io_out_sum_54),
    .io_out_sum_55(accumulation_array_io_out_sum_55),
    .io_out_sum_56(accumulation_array_io_out_sum_56),
    .io_out_sum_57(accumulation_array_io_out_sum_57),
    .io_out_sum_58(accumulation_array_io_out_sum_58),
    .io_out_sum_59(accumulation_array_io_out_sum_59),
    .io_out_sum_60(accumulation_array_io_out_sum_60),
    .io_out_sum_61(accumulation_array_io_out_sum_61),
    .io_out_sum_62(accumulation_array_io_out_sum_62),
    .io_out_sum_63(accumulation_array_io_out_sum_63),
    .io_valid(accumulation_array_io_valid)
  );
  assign io_Data_x_ready = ~activation_buffer_io_isfull; // @[Mini_TPU.scala 85:22]
  assign io_Weight_x_ready = ~weight_buffer_io_isfull; // @[Mini_TPU.scala 80:24]
  assign io_Sum_x_valid = accumulation_array_io_valid; // @[Mini_TPU.scala 90:18]
  assign io_Sum_x_bits_0 = _T_12 ? accumulation_array_io_out_sum_0 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_1 = _T_12 ? accumulation_array_io_out_sum_1 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_2 = _T_12 ? accumulation_array_io_out_sum_2 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_3 = _T_12 ? accumulation_array_io_out_sum_3 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_4 = _T_12 ? accumulation_array_io_out_sum_4 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_5 = _T_12 ? accumulation_array_io_out_sum_5 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_6 = _T_12 ? accumulation_array_io_out_sum_6 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_7 = _T_12 ? accumulation_array_io_out_sum_7 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_8 = _T_12 ? accumulation_array_io_out_sum_8 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_9 = _T_12 ? accumulation_array_io_out_sum_9 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_10 = _T_12 ? accumulation_array_io_out_sum_10 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_11 = _T_12 ? accumulation_array_io_out_sum_11 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_12 = _T_12 ? accumulation_array_io_out_sum_12 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_13 = _T_12 ? accumulation_array_io_out_sum_13 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_14 = _T_12 ? accumulation_array_io_out_sum_14 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_15 = _T_12 ? accumulation_array_io_out_sum_15 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_16 = _T_12 ? accumulation_array_io_out_sum_16 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_17 = _T_12 ? accumulation_array_io_out_sum_17 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_18 = _T_12 ? accumulation_array_io_out_sum_18 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_19 = _T_12 ? accumulation_array_io_out_sum_19 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_20 = _T_12 ? accumulation_array_io_out_sum_20 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_21 = _T_12 ? accumulation_array_io_out_sum_21 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_22 = _T_12 ? accumulation_array_io_out_sum_22 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_23 = _T_12 ? accumulation_array_io_out_sum_23 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_24 = _T_12 ? accumulation_array_io_out_sum_24 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_25 = _T_12 ? accumulation_array_io_out_sum_25 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_26 = _T_12 ? accumulation_array_io_out_sum_26 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_27 = _T_12 ? accumulation_array_io_out_sum_27 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_28 = _T_12 ? accumulation_array_io_out_sum_28 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_29 = _T_12 ? accumulation_array_io_out_sum_29 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_30 = _T_12 ? accumulation_array_io_out_sum_30 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_31 = _T_12 ? accumulation_array_io_out_sum_31 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_32 = _T_12 ? accumulation_array_io_out_sum_32 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_33 = _T_12 ? accumulation_array_io_out_sum_33 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_34 = _T_12 ? accumulation_array_io_out_sum_34 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_35 = _T_12 ? accumulation_array_io_out_sum_35 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_36 = _T_12 ? accumulation_array_io_out_sum_36 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_37 = _T_12 ? accumulation_array_io_out_sum_37 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_38 = _T_12 ? accumulation_array_io_out_sum_38 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_39 = _T_12 ? accumulation_array_io_out_sum_39 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_40 = _T_12 ? accumulation_array_io_out_sum_40 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_41 = _T_12 ? accumulation_array_io_out_sum_41 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_42 = _T_12 ? accumulation_array_io_out_sum_42 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_43 = _T_12 ? accumulation_array_io_out_sum_43 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_44 = _T_12 ? accumulation_array_io_out_sum_44 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_45 = _T_12 ? accumulation_array_io_out_sum_45 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_46 = _T_12 ? accumulation_array_io_out_sum_46 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_47 = _T_12 ? accumulation_array_io_out_sum_47 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_48 = _T_12 ? accumulation_array_io_out_sum_48 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_49 = _T_12 ? accumulation_array_io_out_sum_49 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_50 = _T_12 ? accumulation_array_io_out_sum_50 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_51 = _T_12 ? accumulation_array_io_out_sum_51 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_52 = _T_12 ? accumulation_array_io_out_sum_52 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_53 = _T_12 ? accumulation_array_io_out_sum_53 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_54 = _T_12 ? accumulation_array_io_out_sum_54 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_55 = _T_12 ? accumulation_array_io_out_sum_55 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_56 = _T_12 ? accumulation_array_io_out_sum_56 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_57 = _T_12 ? accumulation_array_io_out_sum_57 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_58 = _T_12 ? accumulation_array_io_out_sum_58 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_59 = _T_12 ? accumulation_array_io_out_sum_59 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_60 = _T_12 ? accumulation_array_io_out_sum_60 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_61 = _T_12 ? accumulation_array_io_out_sum_61 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_62 = _T_12 ? accumulation_array_io_out_sum_62 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign io_Sum_x_bits_63 = _T_12 ? accumulation_array_io_out_sum_63 : 32'h0; // @[Mini_TPU.scala 91:24 92:19 94:19]
  assign activation_buffer_clock = clock;
  assign activation_buffer_reset = reset;
  assign activation_buffer_io_wen = io_Data_x_valid; // @[Mini_TPU.scala 86:28]
  assign activation_buffer_io_ren = 3'h0 == stateReg ? 1'h0 : 3'h1 == stateReg & _GEN_2; // @[Mini_TPU.scala 32:20 27:28]
  assign activation_buffer_io_in_data_x_0 = io_Data_x_bits_0; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_1 = io_Data_x_bits_1; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_2 = io_Data_x_bits_2; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_3 = io_Data_x_bits_3; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_4 = io_Data_x_bits_4; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_5 = io_Data_x_bits_5; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_6 = io_Data_x_bits_6; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_7 = io_Data_x_bits_7; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_8 = io_Data_x_bits_8; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_9 = io_Data_x_bits_9; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_10 = io_Data_x_bits_10; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_11 = io_Data_x_bits_11; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_12 = io_Data_x_bits_12; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_13 = io_Data_x_bits_13; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_14 = io_Data_x_bits_14; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_15 = io_Data_x_bits_15; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_16 = io_Data_x_bits_16; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_17 = io_Data_x_bits_17; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_18 = io_Data_x_bits_18; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_19 = io_Data_x_bits_19; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_20 = io_Data_x_bits_20; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_21 = io_Data_x_bits_21; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_22 = io_Data_x_bits_22; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_23 = io_Data_x_bits_23; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_24 = io_Data_x_bits_24; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_25 = io_Data_x_bits_25; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_26 = io_Data_x_bits_26; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_27 = io_Data_x_bits_27; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_28 = io_Data_x_bits_28; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_29 = io_Data_x_bits_29; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_30 = io_Data_x_bits_30; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_31 = io_Data_x_bits_31; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_32 = io_Data_x_bits_32; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_33 = io_Data_x_bits_33; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_34 = io_Data_x_bits_34; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_35 = io_Data_x_bits_35; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_36 = io_Data_x_bits_36; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_37 = io_Data_x_bits_37; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_38 = io_Data_x_bits_38; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_39 = io_Data_x_bits_39; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_40 = io_Data_x_bits_40; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_41 = io_Data_x_bits_41; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_42 = io_Data_x_bits_42; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_43 = io_Data_x_bits_43; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_44 = io_Data_x_bits_44; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_45 = io_Data_x_bits_45; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_46 = io_Data_x_bits_46; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_47 = io_Data_x_bits_47; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_48 = io_Data_x_bits_48; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_49 = io_Data_x_bits_49; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_50 = io_Data_x_bits_50; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_51 = io_Data_x_bits_51; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_52 = io_Data_x_bits_52; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_53 = io_Data_x_bits_53; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_54 = io_Data_x_bits_54; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_55 = io_Data_x_bits_55; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_56 = io_Data_x_bits_56; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_57 = io_Data_x_bits_57; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_58 = io_Data_x_bits_58; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_59 = io_Data_x_bits_59; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_60 = io_Data_x_bits_60; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_61 = io_Data_x_bits_61; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_62 = io_Data_x_bits_62; // @[Mini_TPU.scala 87:34]
  assign activation_buffer_io_in_data_x_63 = io_Data_x_bits_63; // @[Mini_TPU.scala 87:34]
  assign weight_buffer_clock = clock;
  assign weight_buffer_reset = reset;
  assign weight_buffer_io_wen = io_Weight_x_valid; // @[Mini_TPU.scala 81:24]
  assign weight_buffer_io_ren = 3'h0 == stateReg ? _T_4 : _GEN_21; // @[Mini_TPU.scala 32:20]
  assign weight_buffer_io_in_weight_x_0 = io_Weight_x_bits_0; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_1 = io_Weight_x_bits_1; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_2 = io_Weight_x_bits_2; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_3 = io_Weight_x_bits_3; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_4 = io_Weight_x_bits_4; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_5 = io_Weight_x_bits_5; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_6 = io_Weight_x_bits_6; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_7 = io_Weight_x_bits_7; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_8 = io_Weight_x_bits_8; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_9 = io_Weight_x_bits_9; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_10 = io_Weight_x_bits_10; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_11 = io_Weight_x_bits_11; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_12 = io_Weight_x_bits_12; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_13 = io_Weight_x_bits_13; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_14 = io_Weight_x_bits_14; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_15 = io_Weight_x_bits_15; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_16 = io_Weight_x_bits_16; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_17 = io_Weight_x_bits_17; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_18 = io_Weight_x_bits_18; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_19 = io_Weight_x_bits_19; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_20 = io_Weight_x_bits_20; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_21 = io_Weight_x_bits_21; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_22 = io_Weight_x_bits_22; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_23 = io_Weight_x_bits_23; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_24 = io_Weight_x_bits_24; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_25 = io_Weight_x_bits_25; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_26 = io_Weight_x_bits_26; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_27 = io_Weight_x_bits_27; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_28 = io_Weight_x_bits_28; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_29 = io_Weight_x_bits_29; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_30 = io_Weight_x_bits_30; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_31 = io_Weight_x_bits_31; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_32 = io_Weight_x_bits_32; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_33 = io_Weight_x_bits_33; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_34 = io_Weight_x_bits_34; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_35 = io_Weight_x_bits_35; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_36 = io_Weight_x_bits_36; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_37 = io_Weight_x_bits_37; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_38 = io_Weight_x_bits_38; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_39 = io_Weight_x_bits_39; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_40 = io_Weight_x_bits_40; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_41 = io_Weight_x_bits_41; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_42 = io_Weight_x_bits_42; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_43 = io_Weight_x_bits_43; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_44 = io_Weight_x_bits_44; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_45 = io_Weight_x_bits_45; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_46 = io_Weight_x_bits_46; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_47 = io_Weight_x_bits_47; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_48 = io_Weight_x_bits_48; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_49 = io_Weight_x_bits_49; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_50 = io_Weight_x_bits_50; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_51 = io_Weight_x_bits_51; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_52 = io_Weight_x_bits_52; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_53 = io_Weight_x_bits_53; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_54 = io_Weight_x_bits_54; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_55 = io_Weight_x_bits_55; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_56 = io_Weight_x_bits_56; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_57 = io_Weight_x_bits_57; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_58 = io_Weight_x_bits_58; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_59 = io_Weight_x_bits_59; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_60 = io_Weight_x_bits_60; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_61 = io_Weight_x_bits_61; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_62 = io_Weight_x_bits_62; // @[Mini_TPU.scala 82:32]
  assign weight_buffer_io_in_weight_x_63 = io_Weight_x_bits_63; // @[Mini_TPU.scala 82:32]
  assign systolic_array_clock = clock;
  assign systolic_array_reset = reset;
  assign systolic_array_io_activate_0 = activation_buffer_io_out_activate_0; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_1 = activation_buffer_io_out_activate_1; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_2 = activation_buffer_io_out_activate_2; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_3 = activation_buffer_io_out_activate_3; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_4 = activation_buffer_io_out_activate_4; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_5 = activation_buffer_io_out_activate_5; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_6 = activation_buffer_io_out_activate_6; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_activate_7 = activation_buffer_io_out_activate_7; // @[Mini_TPU.scala 99:30]
  assign systolic_array_io_weight_0 = weight_buffer_io_out_weight_0; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_1 = weight_buffer_io_out_weight_1; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_2 = weight_buffer_io_out_weight_2; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_3 = weight_buffer_io_out_weight_3; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_4 = weight_buffer_io_out_weight_4; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_5 = weight_buffer_io_out_weight_5; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_6 = weight_buffer_io_out_weight_6; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_weight_7 = weight_buffer_io_out_weight_7; // @[Mini_TPU.scala 103:28]
  assign systolic_array_io_flow = activation_buffer_io_out_flow; // @[Mini_TPU.scala 98:26]
  assign systolic_array_io_shift = weight_buffer_io_out_shift; // @[Mini_TPU.scala 102:27]
  assign accumulation_array_clock = clock;
  assign accumulation_array_reset = reset;
  assign accumulation_array_io_in_psum_0 = systolic_array_io_psum_0; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_1 = systolic_array_io_psum_1; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_2 = systolic_array_io_psum_2; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_3 = systolic_array_io_psum_3; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_4 = systolic_array_io_psum_4; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_5 = systolic_array_io_psum_5; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_6 = systolic_array_io_psum_6; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_psum_7 = systolic_array_io_psum_7; // @[Mini_TPU.scala 107:33]
  assign accumulation_array_io_in_valid_0 = systolic_array_io_valid_0; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_1 = systolic_array_io_valid_1; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_2 = systolic_array_io_valid_2; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_3 = systolic_array_io_valid_3; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_4 = systolic_array_io_valid_4; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_5 = systolic_array_io_valid_5; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_6 = systolic_array_io_valid_6; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_valid_7 = systolic_array_io_valid_7; // @[Mini_TPU.scala 106:34]
  assign accumulation_array_io_in_acc = 3'h0 == stateReg ? 1'h0 : _GEN_24; // @[Mini_TPU.scala 32:20 29:32]
  assign accumulation_array_io_in_compute_done = 3'h0 == stateReg ? 1'h0 : _GEN_25; // @[Mini_TPU.scala 32:20 34:45]
  always @(posedge clock) begin
    if (reset) begin // @[Mini_TPU.scala 24:25]
      stateReg <= 3'h0; // @[Mini_TPU.scala 24:25]
    end else if (3'h0 == stateReg) begin // @[Mini_TPU.scala 32:20]
      if (io_Compute & ~activation_buffer_io_isempty & ~weight_buffer_io_isempty) begin // @[Mini_TPU.scala 35:90]
        stateReg <= 3'h1; // @[Mini_TPU.scala 37:18]
      end else begin
        stateReg <= 3'h0; // @[Mini_TPU.scala 39:18]
      end
    end else if (3'h1 == stateReg) begin // @[Mini_TPU.scala 32:20]
      if (weight_buffer_io_isdone) begin // @[Mini_TPU.scala 44:37]
        stateReg <= 3'h2; // @[Mini_TPU.scala 46:18]
      end else begin
        stateReg <= 3'h1; // @[Mini_TPU.scala 48:18]
      end
    end else if (3'h2 == stateReg) begin // @[Mini_TPU.scala 32:20]
      stateReg <= _GEN_5;
    end else begin
      stateReg <= _GEN_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
